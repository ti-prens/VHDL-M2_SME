--*******************************************************************
-- M2 SME 2021/2022
-- BE Synthèse et mise en œuvre des systèmes 
-- Boukah & Jacquet & Ziane 
--*******************************************************************

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
USE ieee.numeric_std.ALL;

--le diviseur dure un cycle d'horloge
entity diviseur is
	generic (
		P : integer := 3 --taille Prescaler
	);
	port (
		Clock, Enable, Reset : in  std_logic;
		Prescaler            : in  std_logic_vector(P-1 downto 0); --prescaler == (PSC + 1) : et doit etre  >=1 
		DivOutput            : out std_logic
	);
end entity diviseur;




architecture rtl of diviseur is
	-- on decl	are les variables d e l'architecture avant le premier begin

	--Prescaler: in std_logic_vector(P-1 downto 0) := 2;

	--signal Prescaler: std_logic_vector(15 downto 0) := x"00ff";
	signal reset_synchrone    : std_logic; -- 1 pour reset synchrone et 0 pour asynchrone
	--signal internal_reset     : std_logic;
	signal sortie_comparateur : std_logic_vector (2 downto 0);
	signal sortie_compteur    : std_logic_vector (P-1 downto 0);
	signal prescaler_value    : std_logic_vector(P-1 downto 0);


	-- declaration des composants
	component comparateur
		--generic ( Q_1 : integer  : = 5);
		generic (
			N : integer
		);
		port (
			valeur_a, valeur_b : in  std_logic_vector (N-1 downto 0);
			sortie_comparaison : out std_logic_vector (2 downto 0)
		-- sortie_comparaison : 100 => a > b ; 010 => a = b ; 001 => a < b
		);
	end component comparateur;


	component compteur is
		generic (
			N : integer
		);
		port (
			clk            : in  std_logic;
			en             : in  std_logic;
			arst_n         : in  std_logic;
			SRst           : in  std_logic;
			counter_output : out std_logic_vector (N-1 downto 0)
		);
	end component compteur;



begin

	prescaler_value <= Prescaler - 1; -- pour avoir 1 coup d'horloge pour chacque prescaler coup d'horloge la comparaison doit se faire sur la valeur precedent le prescler

	U1 : compteur
		generic map (N => P)
		port map(
			clk            => Clock,           --horloge
			en             => Enable,          --enable counting or decounting
			arst_n         => '1',             --reset asynchrone et inverse (1 => pas de reset asynchrone)
			SRst           => reset_synchrone, --reset synchrone
			counter_output => sortie_compteur
		);


	J1 : comparateur -- J1 est une instance du comparateur
		generic map (N => P)
		port map (
			valeur_a           => sortie_compteur,
			valeur_b           => prescaler_value ,
			sortie_comparaison => sortie_comparateur
		); -- remove the 0


	reset_synchrone <= Reset or sortie_comparateur(2);

	-- le comparateur fonctionne en synchrone 
	DivOutput <= sortie_comparateur(1);



end architecture rtl;

--generic ( NomVariable : type  : = "valeur");









