
module nios_mcu (
	clk_clk,
	leds_export,
	reset_reset_n,
	in_freq_anemometre_in_freq_anemometre);	

	input		clk_clk;
	output	[7:0]	leds_export;
	input		reset_reset_n;
	input		in_freq_anemometre_in_freq_anemometre;
endmodule
