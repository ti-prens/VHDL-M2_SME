library IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.ALL;
		  
		  
entity blink is 
	port(
		clk : in bit;
		led : out bit
	);
end entity blink;

architecture rtl of blink is

begin
--

	

end architecture rtl;