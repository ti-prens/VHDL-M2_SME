
module nios_mcu (
	clk_clk,
	in_freq_anemometre_in_freq_anemometre,
	leds_export,
	reset_reset_n);	

	input		clk_clk;
	input		in_freq_anemometre_in_freq_anemometre;
	output	[7:0]	leds_export;
	input		reset_reset_n;
endmodule
