// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition"

// DATE "09/20/2021 11:50:00"

// 
// Device: Altera EP4CE22F17C6 Package FBGA256
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module nios_mcu (
	altera_reserved_tms,
	altera_reserved_tck,
	altera_reserved_tdi,
	altera_reserved_tdo,
	clk_clk,
	leds_export,
	reset_reset_n)/* synthesis synthesis_greybox=1 */;
input 	altera_reserved_tms;
input 	altera_reserved_tck;
input 	altera_reserved_tdi;
output 	altera_reserved_tdo;
input 	clk_clk;
output 	[7:0] leds_export;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[0]~q ;
wire \nios_cpu|cpu|W_alu_result[12]~q ;
wire \nios_cpu|cpu|W_alu_result[15]~q ;
wire \nios_cpu|cpu|W_alu_result[14]~q ;
wire \nios_cpu|cpu|W_alu_result[13]~q ;
wire \nios_cpu|cpu|W_alu_result[11]~q ;
wire \nios_cpu|cpu|W_alu_result[10]~q ;
wire \nios_cpu|cpu|W_alu_result[9]~q ;
wire \nios_cpu|cpu|W_alu_result[8]~q ;
wire \nios_cpu|cpu|W_alu_result[7]~q ;
wire \nios_cpu|cpu|W_alu_result[6]~q ;
wire \nios_cpu|cpu|W_alu_result[5]~q ;
wire \nios_cpu|cpu|W_alu_result[4]~q ;
wire \nios_cpu|cpu|W_alu_result[3]~q ;
wire \nios_cpu|cpu|W_alu_result[2]~q ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[0] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_b[0] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[22] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_b[22] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[23] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_b[23] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[24] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_b[24] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[25] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_b[25] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[26] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_b[26] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[11] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_b[11] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[13] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_b[13] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[16] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_b[16] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[12] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_b[12] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[1] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_b[1] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[3] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_b[3] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[2] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_b[2] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[5] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_b[5] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[4] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_b[4] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[14] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_b[14] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[15] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_b[15] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[18] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_b[18] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[17] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_b[17] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[10] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_b[10] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[9] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_b[9] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[8] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_b[8] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[7] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_b[7] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[6] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_b[6] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[21] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_b[21] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[19] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_b[19] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[20] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_b[20] ;
wire \nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[0]~q ;
wire \nios_cpu|cpu|d_writedata[24]~q ;
wire \nios_cpu|cpu|d_writedata[25]~q ;
wire \nios_cpu|cpu|d_writedata[26]~q ;
wire \nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[1]~q ;
wire \nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[3]~q ;
wire \nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[2]~q ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[27] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_b[27] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[28] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_b[28] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[29] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_b[29] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[30] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_b[30] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_a[31] ;
wire \onchip_ram|the_altsyncram|auto_generated|q_b[31] ;
wire \nios_cpu|cpu|d_writedata[27]~q ;
wire \nios_cpu|cpu|d_writedata[28]~q ;
wire \nios_cpu|cpu|d_writedata[29]~q ;
wire \nios_cpu|cpu|d_writedata[30]~q ;
wire \nios_cpu|cpu|d_writedata[31]~q ;
wire \pio_0|data_out[0]~q ;
wire \pio_0|data_out[1]~q ;
wire \pio_0|data_out[2]~q ;
wire \pio_0|data_out[3]~q ;
wire \pio_0|data_out[4]~q ;
wire \pio_0|data_out[5]~q ;
wire \pio_0|data_out[6]~q ;
wire \pio_0|data_out[7]~q ;
wire \jtag_uart_0|nios_mcu_jtag_uart_0_alt_jtag_atlantic|adapted_tdo~q ;
wire \nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_tck|ir_out[0]~q ;
wire \nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_tck|ir_out[1]~q ;
wire \nios_cpu|cpu|d_writedata[0]~q ;
wire \rst_controller|r_sync_rst~q ;
wire \mm_interconnect_0|router|Equal1~3_combout ;
wire \jtag_uart_0|nios_mcu_jtag_uart_0_alt_jtag_atlantic|rst1~q ;
wire \mm_interconnect_0|pio_0_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \pio_0|always0~0_combout ;
wire \nios_cpu|cpu|d_write~q ;
wire \mm_interconnect_0|nios_cpu_data_master_translator|write_accepted~q ;
wire \mm_interconnect_0|pio_0_s1_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|wait_latency_counter[0]~q ;
wire \nios_cpu|cpu|d_writedata[1]~q ;
wire \nios_cpu|cpu|d_writedata[2]~q ;
wire \nios_cpu|cpu|d_writedata[3]~q ;
wire \nios_cpu|cpu|d_writedata[4]~q ;
wire \nios_cpu|cpu|d_writedata[5]~q ;
wire \nios_cpu|cpu|d_writedata[6]~q ;
wire \nios_cpu|cpu|d_writedata[7]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|read_latency_shift_reg[0]~q ;
wire \nios_cpu|cpu|d_read~q ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg~0_combout ;
wire \mm_interconnect_0|pio_0_s1_agent|m0_write~0_combout ;
wire \mm_interconnect_0|nios_cpu_debug_mem_slave_agent_rsp_fifo|mem[0][73]~q ;
wire \mm_interconnect_0|nios_cpu_debug_mem_slave_agent_rsp_fifo|mem[0][55]~q ;
wire \mm_interconnect_0|nios_cpu_debug_mem_slave_translator|read_latency_shift_reg[0]~q ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg[0]~q ;
wire \mm_interconnect_0|rsp_mux|WideOr1~0_combout ;
wire \mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|read_latency_shift_reg[0]~q ;
wire \mm_interconnect_0|onchip_ram_s2_translator|read_latency_shift_reg[0]~q ;
wire \mm_interconnect_0|rsp_mux|WideOr1~combout ;
wire \mm_interconnect_0|router|Equal3~1_combout ;
wire \mm_interconnect_0|router|src_channel[4]~0_combout ;
wire \mm_interconnect_0|onchip_ram_s2_agent_rsp_fifo|mem_used[1]~q ;
wire \mm_interconnect_0|cmd_mux_002|saved_grant[0]~q ;
wire \nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|the_nios_mcu_nios_cpu_cpu_nios2_ocimem|waitrequest~q ;
wire \mm_interconnect_0|nios_cpu_debug_mem_slave_agent_rsp_fifo|mem_used[1]~q ;
wire \jtag_uart_0|av_waitrequest~q ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_agent_rsp_fifo|mem_used[1]~q ;
wire \mm_interconnect_0|router|Equal2~0_combout ;
wire \avalonslave_0|dRead~q ;
wire \mm_interconnect_0|nios_cpu_data_master_agent|always2~0_combout ;
wire \mm_interconnect_0|avalonslave_0_avalon_slave_0_1_agent|m0_read~0_combout ;
wire \mm_interconnect_0|avalonslave_0_avalon_slave_0_1_agent|m0_read~1_combout ;
wire \avalonslave_0|sReadCountPipelined[0]~32_combout ;
wire \mm_interconnect_0|nios_cpu_data_master_translator|av_waitrequest~2_combout ;
wire \nios_cpu|cpu|F_pc[10]~q ;
wire \nios_cpu|cpu|F_pc[9]~q ;
wire \nios_cpu|cpu|F_pc[8]~q ;
wire \nios_cpu|cpu|F_pc[7]~q ;
wire \nios_cpu|cpu|F_pc[6]~q ;
wire \nios_cpu|cpu|F_pc[5]~q ;
wire \nios_cpu|cpu|F_pc[4]~q ;
wire \nios_cpu|cpu|F_pc[3]~q ;
wire \nios_cpu|cpu|F_pc[2]~q ;
wire \nios_cpu|cpu|F_pc[1]~q ;
wire \nios_cpu|cpu|F_pc[0]~q ;
wire \nios_cpu|cpu|F_pc[13]~q ;
wire \nios_cpu|cpu|F_pc[12]~q ;
wire \nios_cpu|cpu|F_pc[11]~q ;
wire \nios_cpu|cpu|i_read~q ;
wire \mm_interconnect_0|cmd_mux_002|WideOr1~combout ;
wire \avalonslave_0|Equal2~0_combout ;
wire \mm_interconnect_0|nios_cpu_debug_mem_slave_agent|rf_source_valid~1_combout ;
wire \nios_cpu|cpu|hbreak_enabled~q ;
wire \mm_interconnect_0|rsp_mux|WideOr1~1_combout ;
wire \mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[0]~q ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[0]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[0]~q ;
wire \mm_interconnect_0|rsp_demux_002|src0_valid~0_combout ;
wire \mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[0]~q ;
wire \mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[22]~q ;
wire \mm_interconnect_0|onchip_ram_s1_translator|read_latency_shift_reg[0]~q ;
wire \mm_interconnect_0|rsp_demux_002|src1_valid~0_combout ;
wire \mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[23]~q ;
wire \mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[24]~q ;
wire \mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[25]~q ;
wire \mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[26]~q ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~0_combout ;
wire \mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[11]~q ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~1_combout ;
wire \mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[13]~q ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~2_combout ;
wire \mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[16]~q ;
wire \mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[12]~q ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~3_combout ;
wire \mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[1]~q ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~4_combout ;
wire \mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[3]~q ;
wire \mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[2]~q ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~5_combout ;
wire \mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[5]~q ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~6_combout ;
wire \mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[4]~q ;
wire \mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[14]~q ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~7_combout ;
wire \mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[15]~q ;
wire \mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[18]~q ;
wire \mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[17]~q ;
wire \mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[10]~q ;
wire \mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[9]~q ;
wire \mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[8]~q ;
wire \mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[7]~q ;
wire \mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[6]~q ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~8_combout ;
wire \mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[21]~q ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~9_combout ;
wire \mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[19]~q ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~10_combout ;
wire \mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[20]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_data[46]~combout ;
wire \mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[1]~q ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[1]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[1]~q ;
wire \mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[2]~q ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[2]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[2]~q ;
wire \mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[3]~q ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[3]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[3]~q ;
wire \mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[4]~q ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[4]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[4]~q ;
wire \mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[5]~q ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[5]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[5]~q ;
wire \mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[6]~q ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[6]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[6]~q ;
wire \mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[7]~q ;
wire \mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[7]~q ;
wire \mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[7]~q ;
wire \jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_full~q ;
wire \rst_controller|r_early_rst~q ;
wire \mm_interconnect_0|rsp_mux|src_data[8]~1_combout ;
wire \avalonslave_0|ReadData[0]~1_combout ;
wire \jtag_uart_0|read_0~q ;
wire \jtag_uart_0|av_readdata[0]~0_combout ;
wire \nios_cpu|cpu|d_byteenable[0]~q ;
wire \pio_0|readdata[0]~combout ;
wire \jtag_uart_0|av_readdata[9]~combout ;
wire \jtag_uart_0|av_readdata[8]~1_combout ;
wire \nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[22]~q ;
wire \nios_cpu|cpu|d_writedata[22]~q ;
wire \nios_cpu|cpu|d_byteenable[2]~q ;
wire \nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[23]~q ;
wire \nios_cpu|cpu|d_writedata[23]~q ;
wire \nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[24]~q ;
wire \nios_cpu|cpu|d_byteenable[3]~q ;
wire \nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[25]~q ;
wire \nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[26]~q ;
wire \nios_cpu|cpu|d_writedata[11]~q ;
wire \nios_cpu|cpu|d_byteenable[1]~q ;
wire \nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[11]~q ;
wire \nios_cpu|cpu|d_writedata[13]~q ;
wire \nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[13]~q ;
wire \nios_cpu|cpu|d_writedata[16]~q ;
wire \nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[16]~q ;
wire \nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[12]~q ;
wire \nios_cpu|cpu|d_writedata[12]~q ;
wire \nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[5]~q ;
wire \nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[4]~q ;
wire \nios_cpu|cpu|d_writedata[14]~q ;
wire \nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[14]~q ;
wire \nios_cpu|cpu|d_writedata[15]~q ;
wire \nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[15]~q ;
wire \nios_cpu|cpu|d_writedata[18]~q ;
wire \nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[18]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[12]~3_combout ;
wire \mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[27]~q ;
wire \mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[28]~q ;
wire \mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[29]~q ;
wire \mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[30]~q ;
wire \mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[31]~q ;
wire \nios_cpu|cpu|d_writedata[17]~q ;
wire \nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[17]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[11]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[10]~6_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[9]~8_combout ;
wire \nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[10]~q ;
wire \nios_cpu|cpu|d_writedata[10]~q ;
wire \nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[9]~q ;
wire \nios_cpu|cpu|d_writedata[9]~q ;
wire \nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[8]~q ;
wire \nios_cpu|cpu|d_writedata[8]~q ;
wire \nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[7]~q ;
wire \nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[6]~q ;
wire \nios_cpu|cpu|d_writedata[21]~q ;
wire \nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[21]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[15]~10_combout ;
wire \nios_cpu|cpu|d_writedata[19]~q ;
wire \nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[19]~q ;
wire \nios_cpu|cpu|d_writedata[20]~q ;
wire \nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[20]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[14]~12_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[13]~14_combout ;
wire \avalonslave_0|ReadData[1]~3_combout ;
wire \jtag_uart_0|av_readdata[1]~2_combout ;
wire \pio_0|readdata[1]~combout ;
wire \avalonslave_0|ReadData[2]~5_combout ;
wire \jtag_uart_0|av_readdata[2]~3_combout ;
wire \pio_0|readdata[2]~combout ;
wire \avalonslave_0|ReadData[3]~7_combout ;
wire \jtag_uart_0|av_readdata[3]~4_combout ;
wire \pio_0|readdata[3]~combout ;
wire \avalonslave_0|ReadData[4]~9_combout ;
wire \jtag_uart_0|av_readdata[4]~5_combout ;
wire \pio_0|readdata[4]~combout ;
wire \avalonslave_0|ReadData[5]~11_combout ;
wire \jtag_uart_0|av_readdata[5]~6_combout ;
wire \pio_0|readdata[5]~combout ;
wire \avalonslave_0|ReadData[6]~13_combout ;
wire \jtag_uart_0|av_readdata[6]~7_combout ;
wire \pio_0|readdata[6]~combout ;
wire \avalonslave_0|ReadData[7]~15_combout ;
wire \jtag_uart_0|av_readdata[7]~8_combout ;
wire \pio_0|readdata[7]~combout ;
wire \jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ;
wire \jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ;
wire \jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ;
wire \jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ;
wire \jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ;
wire \jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ;
wire \jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~0_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~1_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[38]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[39]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[40]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[41]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[42]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[43]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[44]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[45]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[32]~combout ;
wire \avalonslave_0|ReadData[8]~17_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[16]~16_combout ;
wire \jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ;
wire \jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ;
wire \jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ;
wire \jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ;
wire \jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_full~q ;
wire \jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ;
wire \jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ;
wire \avalonslave_0|ReadData[12]~19_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[20]~18_combout ;
wire \nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[27]~q ;
wire \nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[28]~q ;
wire \nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[29]~q ;
wire \nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[30]~q ;
wire \nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[31]~q ;
wire \avalonslave_0|ReadData[11]~21_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[19]~20_combout ;
wire \avalonslave_0|ReadData[10]~23_combout ;
wire \jtag_uart_0|ac~q ;
wire \mm_interconnect_0|rsp_mux|src_data[18]~22_combout ;
wire \avalonslave_0|ReadData[9]~25_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[17]~24_combout ;
wire \avalonslave_0|ReadData[15]~27_combout ;
wire \jtag_uart_0|rvalid~q ;
wire \mm_interconnect_0|rsp_mux|src_data[23]~combout ;
wire \avalonslave_0|ReadData[14]~29_combout ;
wire \jtag_uart_0|woverflow~q ;
wire \mm_interconnect_0|rsp_mux|src_data[22]~27_combout ;
wire \avalonslave_0|ReadData[13]~31_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[21]~29_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~2_combout ;
wire \avalonslave_0|ReadData[16]~33_combout ;
wire \mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[24]~q ;
wire \mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[31]~q ;
wire \mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[30]~q ;
wire \mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[29]~q ;
wire \mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[28]~q ;
wire \mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[27]~q ;
wire \mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[26]~q ;
wire \mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[25]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~3_combout ;
wire \avalonslave_0|ReadData[20]~35_combout ;
wire \avalonslave_0|ReadData[19]~37_combout ;
wire \avalonslave_0|ReadData[18]~39_combout ;
wire \avalonslave_0|ReadData[17]~41_combout ;
wire \avalonslave_0|ReadData[23]~43_combout ;
wire \avalonslave_0|ReadData[22]~45_combout ;
wire \avalonslave_0|ReadData[21]~47_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~4_combout ;
wire \avalonslave_0|ReadData[24]~49_combout ;
wire \avalonslave_0|ReadData[31]~51_combout ;
wire \avalonslave_0|ReadData[30]~53_combout ;
wire \avalonslave_0|ReadData[29]~55_combout ;
wire \avalonslave_0|ReadData[28]~57_combout ;
wire \avalonslave_0|ReadData[27]~59_combout ;
wire \avalonslave_0|ReadData[26]~61_combout ;
wire \avalonslave_0|ReadData[25]~63_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~5_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[34]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~6_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~7_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[35]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~8_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~9_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~10_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[33]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~11_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~12_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~13_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~14_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~15_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~16_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~17_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~18_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~19_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~20_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~21_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~22_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~23_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~24_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~25_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~26_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~27_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~28_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~29_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~30_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~31_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~32_combout ;
wire \rst_controller|alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain[1]~0_combout ;
wire \~GND~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~8_combout ;
wire \auto_hub|~GND~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ;
wire \clk_clk~input_o ;
wire \reset_reset_n~input_o ;
wire \altera_reserved_tms~input_o ;
wire \altera_reserved_tck~input_o ;
wire \altera_reserved_tdi~input_o ;
wire \altera_internal_jtag~TCKUTAP ;
wire \altera_internal_jtag~TMSUTAP ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ;
wire \altera_internal_jtag~TDIUTAP ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~14_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~16_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~15_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~10 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~13 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~14_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~15 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~16_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~17 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~18_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~20_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~16_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~17_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~18_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~19_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~20_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~25_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~26_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~23_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~24_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~21_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~22_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~23_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~19_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~22_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~12 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~14 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~15_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~17_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~14_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~16_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~17_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~19_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~15_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~18_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ;
wire \altera_internal_jtag~TDO ;


nios_mcu_nios_mcu_nios_cpu nios_cpu(
	.sr_0(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[0]~q ),
	.W_alu_result_12(\nios_cpu|cpu|W_alu_result[12]~q ),
	.W_alu_result_15(\nios_cpu|cpu|W_alu_result[15]~q ),
	.W_alu_result_14(\nios_cpu|cpu|W_alu_result[14]~q ),
	.W_alu_result_13(\nios_cpu|cpu|W_alu_result[13]~q ),
	.W_alu_result_11(\nios_cpu|cpu|W_alu_result[11]~q ),
	.W_alu_result_10(\nios_cpu|cpu|W_alu_result[10]~q ),
	.W_alu_result_9(\nios_cpu|cpu|W_alu_result[9]~q ),
	.W_alu_result_8(\nios_cpu|cpu|W_alu_result[8]~q ),
	.W_alu_result_7(\nios_cpu|cpu|W_alu_result[7]~q ),
	.W_alu_result_6(\nios_cpu|cpu|W_alu_result[6]~q ),
	.W_alu_result_5(\nios_cpu|cpu|W_alu_result[5]~q ),
	.W_alu_result_4(\nios_cpu|cpu|W_alu_result[4]~q ),
	.W_alu_result_3(\nios_cpu|cpu|W_alu_result[3]~q ),
	.W_alu_result_2(\nios_cpu|cpu|W_alu_result[2]~q ),
	.q_a_0(\onchip_ram|the_altsyncram|auto_generated|q_a[0] ),
	.q_b_0(\onchip_ram|the_altsyncram|auto_generated|q_b[0] ),
	.q_a_22(\onchip_ram|the_altsyncram|auto_generated|q_a[22] ),
	.q_a_23(\onchip_ram|the_altsyncram|auto_generated|q_a[23] ),
	.q_a_24(\onchip_ram|the_altsyncram|auto_generated|q_a[24] ),
	.q_b_24(\onchip_ram|the_altsyncram|auto_generated|q_b[24] ),
	.q_a_25(\onchip_ram|the_altsyncram|auto_generated|q_a[25] ),
	.q_b_25(\onchip_ram|the_altsyncram|auto_generated|q_b[25] ),
	.q_a_26(\onchip_ram|the_altsyncram|auto_generated|q_a[26] ),
	.q_b_26(\onchip_ram|the_altsyncram|auto_generated|q_b[26] ),
	.q_a_12(\onchip_ram|the_altsyncram|auto_generated|q_a[12] ),
	.q_b_1(\onchip_ram|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_3(\onchip_ram|the_altsyncram|auto_generated|q_b[3] ),
	.q_a_2(\onchip_ram|the_altsyncram|auto_generated|q_a[2] ),
	.q_b_2(\onchip_ram|the_altsyncram|auto_generated|q_b[2] ),
	.q_b_5(\onchip_ram|the_altsyncram|auto_generated|q_b[5] ),
	.q_b_4(\onchip_ram|the_altsyncram|auto_generated|q_b[4] ),
	.q_a_14(\onchip_ram|the_altsyncram|auto_generated|q_a[14] ),
	.q_a_18(\onchip_ram|the_altsyncram|auto_generated|q_a[18] ),
	.q_a_17(\onchip_ram|the_altsyncram|auto_generated|q_a[17] ),
	.q_a_10(\onchip_ram|the_altsyncram|auto_generated|q_a[10] ),
	.q_a_9(\onchip_ram|the_altsyncram|auto_generated|q_a[9] ),
	.q_a_8(\onchip_ram|the_altsyncram|auto_generated|q_a[8] ),
	.q_a_7(\onchip_ram|the_altsyncram|auto_generated|q_a[7] ),
	.q_b_7(\onchip_ram|the_altsyncram|auto_generated|q_b[7] ),
	.q_a_6(\onchip_ram|the_altsyncram|auto_generated|q_a[6] ),
	.q_b_6(\onchip_ram|the_altsyncram|auto_generated|q_b[6] ),
	.readdata_0(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[0]~q ),
	.d_writedata_24(\nios_cpu|cpu|d_writedata[24]~q ),
	.d_writedata_25(\nios_cpu|cpu|d_writedata[25]~q ),
	.d_writedata_26(\nios_cpu|cpu|d_writedata[26]~q ),
	.readdata_1(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[1]~q ),
	.readdata_3(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[3]~q ),
	.readdata_2(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[2]~q ),
	.q_a_27(\onchip_ram|the_altsyncram|auto_generated|q_a[27] ),
	.q_b_27(\onchip_ram|the_altsyncram|auto_generated|q_b[27] ),
	.q_a_28(\onchip_ram|the_altsyncram|auto_generated|q_a[28] ),
	.q_b_28(\onchip_ram|the_altsyncram|auto_generated|q_b[28] ),
	.q_a_29(\onchip_ram|the_altsyncram|auto_generated|q_a[29] ),
	.q_b_29(\onchip_ram|the_altsyncram|auto_generated|q_b[29] ),
	.q_a_30(\onchip_ram|the_altsyncram|auto_generated|q_a[30] ),
	.q_b_30(\onchip_ram|the_altsyncram|auto_generated|q_b[30] ),
	.q_a_31(\onchip_ram|the_altsyncram|auto_generated|q_a[31] ),
	.q_b_31(\onchip_ram|the_altsyncram|auto_generated|q_b[31] ),
	.d_writedata_27(\nios_cpu|cpu|d_writedata[27]~q ),
	.d_writedata_28(\nios_cpu|cpu|d_writedata[28]~q ),
	.d_writedata_29(\nios_cpu|cpu|d_writedata[29]~q ),
	.d_writedata_30(\nios_cpu|cpu|d_writedata[30]~q ),
	.d_writedata_31(\nios_cpu|cpu|d_writedata[31]~q ),
	.ir_out_0(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_tck|ir_out[0]~q ),
	.ir_out_1(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_tck|ir_out[1]~q ),
	.d_writedata_0(\nios_cpu|cpu|d_writedata[0]~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.d_write(\nios_cpu|cpu|d_write~q ),
	.d_writedata_1(\nios_cpu|cpu|d_writedata[1]~q ),
	.d_writedata_2(\nios_cpu|cpu|d_writedata[2]~q ),
	.d_writedata_3(\nios_cpu|cpu|d_writedata[3]~q ),
	.d_writedata_4(\nios_cpu|cpu|d_writedata[4]~q ),
	.d_writedata_5(\nios_cpu|cpu|d_writedata[5]~q ),
	.d_writedata_6(\nios_cpu|cpu|d_writedata[6]~q ),
	.d_writedata_7(\nios_cpu|cpu|d_writedata[7]~q ),
	.read_latency_shift_reg_0(\mm_interconnect_0|pio_0_s1_translator|read_latency_shift_reg[0]~q ),
	.d_read(\nios_cpu|cpu|d_read~q ),
	.m0_write(\mm_interconnect_0|pio_0_s1_agent|m0_write~0_combout ),
	.mem_73_0(\mm_interconnect_0|nios_cpu_debug_mem_slave_agent_rsp_fifo|mem[0][73]~q ),
	.mem_55_0(\mm_interconnect_0|nios_cpu_debug_mem_slave_agent_rsp_fifo|mem[0][55]~q ),
	.read_latency_shift_reg_01(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_02(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg[0]~q ),
	.WideOr1(\mm_interconnect_0|rsp_mux|WideOr1~0_combout ),
	.read_latency_shift_reg_03(\mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_04(\mm_interconnect_0|onchip_ram_s2_translator|read_latency_shift_reg[0]~q ),
	.WideOr11(\mm_interconnect_0|rsp_mux|WideOr1~combout ),
	.saved_grant_0(\mm_interconnect_0|cmd_mux_002|saved_grant[0]~q ),
	.debug_mem_slave_waitrequest(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|the_nios_mcu_nios_cpu_cpu_nios2_ocimem|waitrequest~q ),
	.mem_used_1(\mm_interconnect_0|nios_cpu_debug_mem_slave_agent_rsp_fifo|mem_used[1]~q ),
	.av_waitrequest(\mm_interconnect_0|nios_cpu_data_master_translator|av_waitrequest~2_combout ),
	.F_pc_10(\nios_cpu|cpu|F_pc[10]~q ),
	.F_pc_9(\nios_cpu|cpu|F_pc[9]~q ),
	.F_pc_8(\nios_cpu|cpu|F_pc[8]~q ),
	.F_pc_7(\nios_cpu|cpu|F_pc[7]~q ),
	.F_pc_6(\nios_cpu|cpu|F_pc[6]~q ),
	.F_pc_5(\nios_cpu|cpu|F_pc[5]~q ),
	.F_pc_4(\nios_cpu|cpu|F_pc[4]~q ),
	.F_pc_3(\nios_cpu|cpu|F_pc[3]~q ),
	.F_pc_2(\nios_cpu|cpu|F_pc[2]~q ),
	.F_pc_1(\nios_cpu|cpu|F_pc[1]~q ),
	.F_pc_0(\nios_cpu|cpu|F_pc[0]~q ),
	.F_pc_13(\nios_cpu|cpu|F_pc[13]~q ),
	.F_pc_12(\nios_cpu|cpu|F_pc[12]~q ),
	.F_pc_11(\nios_cpu|cpu|F_pc[11]~q ),
	.i_read(\nios_cpu|cpu|i_read~q ),
	.WideOr12(\mm_interconnect_0|cmd_mux_002|WideOr1~combout ),
	.rf_source_valid(\mm_interconnect_0|nios_cpu_debug_mem_slave_agent|rf_source_valid~1_combout ),
	.hbreak_enabled(\nios_cpu|cpu|hbreak_enabled~q ),
	.WideOr13(\mm_interconnect_0|rsp_mux|WideOr1~1_combout ),
	.av_readdata_pre_0(\mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_01(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_02(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[0]~q ),
	.src0_valid(\mm_interconnect_0|rsp_demux_002|src0_valid~0_combout ),
	.av_readdata_pre_03(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_22(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[22]~q ),
	.read_latency_shift_reg_05(\mm_interconnect_0|onchip_ram_s1_translator|read_latency_shift_reg[0]~q ),
	.src1_valid(\mm_interconnect_0|rsp_demux_002|src1_valid~0_combout ),
	.av_readdata_pre_23(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[23]~q ),
	.av_readdata_pre_24(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[24]~q ),
	.av_readdata_pre_25(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[25]~q ),
	.av_readdata_pre_26(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[26]~q ),
	.src_payload(\mm_interconnect_0|rsp_mux_001|src_payload~0_combout ),
	.av_readdata_pre_11(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[11]~q ),
	.src_payload1(\mm_interconnect_0|rsp_mux_001|src_payload~1_combout ),
	.av_readdata_pre_13(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[13]~q ),
	.src_payload2(\mm_interconnect_0|rsp_mux_001|src_payload~2_combout ),
	.av_readdata_pre_16(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[16]~q ),
	.av_readdata_pre_12(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[12]~q ),
	.src_payload3(\mm_interconnect_0|rsp_mux_001|src_payload~3_combout ),
	.av_readdata_pre_1(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[1]~q ),
	.src_payload4(\mm_interconnect_0|rsp_mux_001|src_payload~4_combout ),
	.av_readdata_pre_3(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_2(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[2]~q ),
	.src_payload5(\mm_interconnect_0|rsp_mux_001|src_payload~5_combout ),
	.av_readdata_pre_5(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[5]~q ),
	.src_payload6(\mm_interconnect_0|rsp_mux_001|src_payload~6_combout ),
	.av_readdata_pre_4(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_14(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[14]~q ),
	.src_payload7(\mm_interconnect_0|rsp_mux_001|src_payload~7_combout ),
	.av_readdata_pre_15(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_18(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[18]~q ),
	.av_readdata_pre_17(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[17]~q ),
	.av_readdata_pre_10(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_9(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_8(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_7(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_6(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[6]~q ),
	.src_payload8(\mm_interconnect_0|rsp_mux_001|src_payload~8_combout ),
	.av_readdata_pre_21(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[21]~q ),
	.src_payload9(\mm_interconnect_0|rsp_mux_001|src_payload~9_combout ),
	.av_readdata_pre_19(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[19]~q ),
	.src_payload10(\mm_interconnect_0|rsp_mux_001|src_payload~10_combout ),
	.av_readdata_pre_20(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[20]~q ),
	.src_data_46(\mm_interconnect_0|cmd_mux_002|src_data[46]~combout ),
	.av_readdata_pre_110(\mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_111(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_112(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_27(\mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_28(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_29(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_31(\mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_32(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_33(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_41(\mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_42(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_43(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_51(\mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_52(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_53(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_61(\mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_62(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_63(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_71(\mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_72(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_73(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[7]~q ),
	.r_early_rst(\rst_controller|r_early_rst~q ),
	.src_data_8(\mm_interconnect_0|rsp_mux|src_data[8]~1_combout ),
	.d_byteenable_0(\nios_cpu|cpu|d_byteenable[0]~q ),
	.av_readdata_9(\jtag_uart_0|av_readdata[9]~combout ),
	.av_readdata_8(\jtag_uart_0|av_readdata[8]~1_combout ),
	.readdata_22(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[22]~q ),
	.d_writedata_22(\nios_cpu|cpu|d_writedata[22]~q ),
	.d_byteenable_2(\nios_cpu|cpu|d_byteenable[2]~q ),
	.readdata_23(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[23]~q ),
	.d_writedata_23(\nios_cpu|cpu|d_writedata[23]~q ),
	.readdata_24(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[24]~q ),
	.d_byteenable_3(\nios_cpu|cpu|d_byteenable[3]~q ),
	.readdata_25(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[25]~q ),
	.readdata_26(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[26]~q ),
	.d_writedata_11(\nios_cpu|cpu|d_writedata[11]~q ),
	.d_byteenable_1(\nios_cpu|cpu|d_byteenable[1]~q ),
	.readdata_11(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[11]~q ),
	.d_writedata_13(\nios_cpu|cpu|d_writedata[13]~q ),
	.readdata_13(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[13]~q ),
	.d_writedata_16(\nios_cpu|cpu|d_writedata[16]~q ),
	.readdata_16(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[16]~q ),
	.readdata_12(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[12]~q ),
	.d_writedata_12(\nios_cpu|cpu|d_writedata[12]~q ),
	.readdata_5(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[5]~q ),
	.readdata_4(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[4]~q ),
	.d_writedata_14(\nios_cpu|cpu|d_writedata[14]~q ),
	.readdata_14(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[14]~q ),
	.d_writedata_15(\nios_cpu|cpu|d_writedata[15]~q ),
	.readdata_15(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[15]~q ),
	.d_writedata_18(\nios_cpu|cpu|d_writedata[18]~q ),
	.readdata_18(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[18]~q ),
	.src_data_12(\mm_interconnect_0|rsp_mux|src_data[12]~3_combout ),
	.av_readdata_pre_271(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[27]~q ),
	.av_readdata_pre_281(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[28]~q ),
	.av_readdata_pre_291(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[29]~q ),
	.av_readdata_pre_30(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[30]~q ),
	.av_readdata_pre_311(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[31]~q ),
	.d_writedata_17(\nios_cpu|cpu|d_writedata[17]~q ),
	.readdata_17(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[17]~q ),
	.src_data_11(\mm_interconnect_0|rsp_mux|src_data[11]~combout ),
	.src_data_10(\mm_interconnect_0|rsp_mux|src_data[10]~6_combout ),
	.src_data_9(\mm_interconnect_0|rsp_mux|src_data[9]~8_combout ),
	.readdata_10(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[10]~q ),
	.d_writedata_10(\nios_cpu|cpu|d_writedata[10]~q ),
	.readdata_9(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[9]~q ),
	.d_writedata_9(\nios_cpu|cpu|d_writedata[9]~q ),
	.readdata_8(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[8]~q ),
	.d_writedata_8(\nios_cpu|cpu|d_writedata[8]~q ),
	.readdata_7(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[7]~q ),
	.readdata_6(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[6]~q ),
	.d_writedata_21(\nios_cpu|cpu|d_writedata[21]~q ),
	.readdata_21(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[21]~q ),
	.src_data_15(\mm_interconnect_0|rsp_mux|src_data[15]~10_combout ),
	.d_writedata_19(\nios_cpu|cpu|d_writedata[19]~q ),
	.readdata_19(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[19]~q ),
	.d_writedata_20(\nios_cpu|cpu|d_writedata[20]~q ),
	.readdata_20(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[20]~q ),
	.src_data_14(\mm_interconnect_0|rsp_mux|src_data[14]~12_combout ),
	.src_data_13(\mm_interconnect_0|rsp_mux|src_data[13]~14_combout ),
	.src_payload11(\mm_interconnect_0|cmd_mux_002|src_payload~0_combout ),
	.src_payload12(\mm_interconnect_0|cmd_mux_002|src_payload~1_combout ),
	.src_data_38(\mm_interconnect_0|cmd_mux_002|src_data[38]~combout ),
	.src_data_39(\mm_interconnect_0|cmd_mux_002|src_data[39]~combout ),
	.src_data_40(\mm_interconnect_0|cmd_mux_002|src_data[40]~combout ),
	.src_data_41(\mm_interconnect_0|cmd_mux_002|src_data[41]~combout ),
	.src_data_42(\mm_interconnect_0|cmd_mux_002|src_data[42]~combout ),
	.src_data_43(\mm_interconnect_0|cmd_mux_002|src_data[43]~combout ),
	.src_data_44(\mm_interconnect_0|cmd_mux_002|src_data[44]~combout ),
	.src_data_45(\mm_interconnect_0|cmd_mux_002|src_data[45]~combout ),
	.src_data_32(\mm_interconnect_0|cmd_mux_002|src_data[32]~combout ),
	.src_data_16(\mm_interconnect_0|rsp_mux|src_data[16]~16_combout ),
	.src_data_20(\mm_interconnect_0|rsp_mux|src_data[20]~18_combout ),
	.readdata_27(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[27]~q ),
	.readdata_28(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[28]~q ),
	.readdata_29(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[29]~q ),
	.readdata_30(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[30]~q ),
	.readdata_31(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[31]~q ),
	.src_data_19(\mm_interconnect_0|rsp_mux|src_data[19]~20_combout ),
	.src_data_18(\mm_interconnect_0|rsp_mux|src_data[18]~22_combout ),
	.src_data_17(\mm_interconnect_0|rsp_mux|src_data[17]~24_combout ),
	.src_data_23(\mm_interconnect_0|rsp_mux|src_data[23]~combout ),
	.src_data_22(\mm_interconnect_0|rsp_mux|src_data[22]~27_combout ),
	.src_data_21(\mm_interconnect_0|rsp_mux|src_data[21]~29_combout ),
	.src_payload13(\mm_interconnect_0|cmd_mux_002|src_payload~2_combout ),
	.av_readdata_pre_241(\mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[24]~q ),
	.av_readdata_pre_312(\mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[31]~q ),
	.av_readdata_pre_301(\mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[30]~q ),
	.av_readdata_pre_292(\mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[29]~q ),
	.av_readdata_pre_282(\mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[28]~q ),
	.av_readdata_pre_272(\mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[27]~q ),
	.av_readdata_pre_261(\mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[26]~q ),
	.av_readdata_pre_251(\mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[25]~q ),
	.src_payload14(\mm_interconnect_0|cmd_mux_002|src_payload~3_combout ),
	.src_payload15(\mm_interconnect_0|cmd_mux_002|src_payload~4_combout ),
	.src_payload16(\mm_interconnect_0|cmd_mux_002|src_payload~5_combout ),
	.src_data_34(\mm_interconnect_0|cmd_mux_002|src_data[34]~combout ),
	.src_payload17(\mm_interconnect_0|cmd_mux_002|src_payload~6_combout ),
	.src_payload18(\mm_interconnect_0|cmd_mux_002|src_payload~7_combout ),
	.src_data_35(\mm_interconnect_0|cmd_mux_002|src_data[35]~combout ),
	.src_payload19(\mm_interconnect_0|cmd_mux_002|src_payload~8_combout ),
	.src_payload20(\mm_interconnect_0|cmd_mux_002|src_payload~9_combout ),
	.src_payload21(\mm_interconnect_0|cmd_mux_002|src_payload~10_combout ),
	.src_data_33(\mm_interconnect_0|cmd_mux_002|src_data[33]~combout ),
	.src_payload22(\mm_interconnect_0|cmd_mux_002|src_payload~11_combout ),
	.src_payload23(\mm_interconnect_0|cmd_mux_002|src_payload~12_combout ),
	.src_payload24(\mm_interconnect_0|cmd_mux_002|src_payload~13_combout ),
	.src_payload25(\mm_interconnect_0|cmd_mux_002|src_payload~14_combout ),
	.src_payload26(\mm_interconnect_0|cmd_mux_002|src_payload~15_combout ),
	.src_payload27(\mm_interconnect_0|cmd_mux_002|src_payload~16_combout ),
	.src_payload28(\mm_interconnect_0|cmd_mux_002|src_payload~17_combout ),
	.src_payload29(\mm_interconnect_0|cmd_mux_002|src_payload~18_combout ),
	.src_payload30(\mm_interconnect_0|cmd_mux_002|src_payload~19_combout ),
	.src_payload31(\mm_interconnect_0|cmd_mux_002|src_payload~20_combout ),
	.src_payload32(\mm_interconnect_0|cmd_mux_002|src_payload~21_combout ),
	.src_payload33(\mm_interconnect_0|cmd_mux_002|src_payload~22_combout ),
	.src_payload34(\mm_interconnect_0|cmd_mux_002|src_payload~23_combout ),
	.src_payload35(\mm_interconnect_0|cmd_mux_002|src_payload~24_combout ),
	.src_payload36(\mm_interconnect_0|cmd_mux_002|src_payload~25_combout ),
	.src_payload37(\mm_interconnect_0|cmd_mux_002|src_payload~26_combout ),
	.src_payload38(\mm_interconnect_0|cmd_mux_002|src_payload~27_combout ),
	.src_payload39(\mm_interconnect_0|cmd_mux_002|src_payload~28_combout ),
	.src_payload40(\mm_interconnect_0|cmd_mux_002|src_payload~29_combout ),
	.src_payload41(\mm_interconnect_0|cmd_mux_002|src_payload~30_combout ),
	.src_payload42(\mm_interconnect_0|cmd_mux_002|src_payload~31_combout ),
	.src_payload43(\mm_interconnect_0|cmd_mux_002|src_payload~32_combout ),
	.altera_internal_jtag(\altera_internal_jtag~TCKUTAP ),
	.altera_internal_jtag1(\altera_internal_jtag~TDIUTAP ),
	.state_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.state_4(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.virtual_ir_scan_reg(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.state_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.state_8(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.splitter_nodes_receive_1_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3]~q ),
	.irf_reg_0_2(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ),
	.irf_reg_1_2(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ),
	.clk_clk(\clk_clk~input_o ));

nios_mcu_nios_mcu_jtag_uart_0 jtag_uart_0(
	.W_alu_result_2(\nios_cpu|cpu|W_alu_result[2]~q ),
	.adapted_tdo(\jtag_uart_0|nios_mcu_jtag_uart_0_alt_jtag_atlantic|adapted_tdo~q ),
	.d_writedata_0(\nios_cpu|cpu|d_writedata[0]~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.rst1(\jtag_uart_0|nios_mcu_jtag_uart_0_alt_jtag_atlantic|rst1~q ),
	.d_writedata_1(\nios_cpu|cpu|d_writedata[1]~q ),
	.d_writedata_2(\nios_cpu|cpu|d_writedata[2]~q ),
	.d_writedata_3(\nios_cpu|cpu|d_writedata[3]~q ),
	.d_writedata_4(\nios_cpu|cpu|d_writedata[4]~q ),
	.d_writedata_5(\nios_cpu|cpu|d_writedata[5]~q ),
	.d_writedata_6(\nios_cpu|cpu|d_writedata[6]~q ),
	.d_writedata_7(\nios_cpu|cpu|d_writedata[7]~q ),
	.read_latency_shift_reg(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg~0_combout ),
	.m0_write(\mm_interconnect_0|pio_0_s1_agent|m0_write~0_combout ),
	.Equal3(\mm_interconnect_0|router|Equal3~1_combout ),
	.av_waitrequest1(\jtag_uart_0|av_waitrequest~q ),
	.mem_used_1(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_agent_rsp_fifo|mem_used[1]~q ),
	.always2(\mm_interconnect_0|nios_cpu_data_master_agent|always2~0_combout ),
	.b_full(\jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.read_01(\jtag_uart_0|read_0~q ),
	.av_readdata_0(\jtag_uart_0|av_readdata[0]~0_combout ),
	.av_readdata_9(\jtag_uart_0|av_readdata[9]~combout ),
	.av_readdata_8(\jtag_uart_0|av_readdata[8]~1_combout ),
	.d_writedata_10(\nios_cpu|cpu|d_writedata[10]~q ),
	.av_readdata_1(\jtag_uart_0|av_readdata[1]~2_combout ),
	.av_readdata_2(\jtag_uart_0|av_readdata[2]~3_combout ),
	.av_readdata_3(\jtag_uart_0|av_readdata[3]~4_combout ),
	.av_readdata_4(\jtag_uart_0|av_readdata[4]~5_combout ),
	.av_readdata_5(\jtag_uart_0|av_readdata[5]~6_combout ),
	.av_readdata_6(\jtag_uart_0|av_readdata[6]~7_combout ),
	.av_readdata_7(\jtag_uart_0|av_readdata[7]~8_combout ),
	.b_non_empty(\jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.counter_reg_bit_5(\jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.counter_reg_bit_4(\jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.counter_reg_bit_2(\jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.counter_reg_bit_31(\jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.counter_reg_bit_01(\jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.counter_reg_bit_21(\jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.counter_reg_bit_11(\jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.b_full1(\jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.counter_reg_bit_51(\jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.counter_reg_bit_41(\jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.ac1(\jtag_uart_0|ac~q ),
	.rvalid1(\jtag_uart_0|rvalid~q ),
	.woverflow1(\jtag_uart_0|woverflow~q ),
	.altera_internal_jtag(\altera_internal_jtag~TCKUTAP ),
	.altera_internal_jtag1(\altera_internal_jtag~TDIUTAP ),
	.state_4(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.splitter_nodes_receive_0_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.virtual_ir_scan_reg(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.clr_reg(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.state_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.state_8(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.irf_reg_0_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.clk_clk(\clk_clk~input_o ));

nios_mcu_AvalonSlave avalonslave_0(
	.W_alu_result_3(\nios_cpu|cpu|W_alu_result[3]~q ),
	.W_alu_result_2(\nios_cpu|cpu|W_alu_result[2]~q ),
	.d_writedata_24(\nios_cpu|cpu|d_writedata[24]~q ),
	.d_writedata_25(\nios_cpu|cpu|d_writedata[25]~q ),
	.d_writedata_26(\nios_cpu|cpu|d_writedata[26]~q ),
	.d_writedata_27(\nios_cpu|cpu|d_writedata[27]~q ),
	.d_writedata_28(\nios_cpu|cpu|d_writedata[28]~q ),
	.d_writedata_29(\nios_cpu|cpu|d_writedata[29]~q ),
	.d_writedata_30(\nios_cpu|cpu|d_writedata[30]~q ),
	.d_writedata_31(\nios_cpu|cpu|d_writedata[31]~q ),
	.d_writedata_0(\nios_cpu|cpu|d_writedata[0]~q ),
	.d_writedata_1(\nios_cpu|cpu|d_writedata[1]~q ),
	.d_writedata_2(\nios_cpu|cpu|d_writedata[2]~q ),
	.d_writedata_3(\nios_cpu|cpu|d_writedata[3]~q ),
	.d_writedata_4(\nios_cpu|cpu|d_writedata[4]~q ),
	.d_writedata_5(\nios_cpu|cpu|d_writedata[5]~q ),
	.d_writedata_6(\nios_cpu|cpu|d_writedata[6]~q ),
	.d_writedata_7(\nios_cpu|cpu|d_writedata[7]~q ),
	.m0_write(\mm_interconnect_0|pio_0_s1_agent|m0_write~0_combout ),
	.Equal2(\mm_interconnect_0|router|Equal2~0_combout ),
	.dRead1(\avalonslave_0|dRead~q ),
	.m0_read(\mm_interconnect_0|avalonslave_0_avalon_slave_0_1_agent|m0_read~0_combout ),
	.Read(\mm_interconnect_0|avalonslave_0_avalon_slave_0_1_agent|m0_read~1_combout ),
	.sReadCountPipelined_0(\avalonslave_0|sReadCountPipelined[0]~32_combout ),
	.Equal21(\avalonslave_0|Equal2~0_combout ),
	.ReadData_0(\avalonslave_0|ReadData[0]~1_combout ),
	.d_byteenable_0(\nios_cpu|cpu|d_byteenable[0]~q ),
	.d_writedata_22(\nios_cpu|cpu|d_writedata[22]~q ),
	.d_byteenable_2(\nios_cpu|cpu|d_byteenable[2]~q ),
	.d_writedata_23(\nios_cpu|cpu|d_writedata[23]~q ),
	.d_byteenable_3(\nios_cpu|cpu|d_byteenable[3]~q ),
	.d_writedata_11(\nios_cpu|cpu|d_writedata[11]~q ),
	.d_byteenable_1(\nios_cpu|cpu|d_byteenable[1]~q ),
	.d_writedata_13(\nios_cpu|cpu|d_writedata[13]~q ),
	.d_writedata_16(\nios_cpu|cpu|d_writedata[16]~q ),
	.d_writedata_12(\nios_cpu|cpu|d_writedata[12]~q ),
	.d_writedata_14(\nios_cpu|cpu|d_writedata[14]~q ),
	.d_writedata_15(\nios_cpu|cpu|d_writedata[15]~q ),
	.d_writedata_18(\nios_cpu|cpu|d_writedata[18]~q ),
	.d_writedata_17(\nios_cpu|cpu|d_writedata[17]~q ),
	.d_writedata_10(\nios_cpu|cpu|d_writedata[10]~q ),
	.d_writedata_9(\nios_cpu|cpu|d_writedata[9]~q ),
	.d_writedata_8(\nios_cpu|cpu|d_writedata[8]~q ),
	.d_writedata_21(\nios_cpu|cpu|d_writedata[21]~q ),
	.d_writedata_19(\nios_cpu|cpu|d_writedata[19]~q ),
	.d_writedata_20(\nios_cpu|cpu|d_writedata[20]~q ),
	.ReadData_1(\avalonslave_0|ReadData[1]~3_combout ),
	.ReadData_2(\avalonslave_0|ReadData[2]~5_combout ),
	.ReadData_3(\avalonslave_0|ReadData[3]~7_combout ),
	.ReadData_4(\avalonslave_0|ReadData[4]~9_combout ),
	.ReadData_5(\avalonslave_0|ReadData[5]~11_combout ),
	.ReadData_6(\avalonslave_0|ReadData[6]~13_combout ),
	.ReadData_7(\avalonslave_0|ReadData[7]~15_combout ),
	.ReadData_8(\avalonslave_0|ReadData[8]~17_combout ),
	.ReadData_12(\avalonslave_0|ReadData[12]~19_combout ),
	.ReadData_11(\avalonslave_0|ReadData[11]~21_combout ),
	.ReadData_10(\avalonslave_0|ReadData[10]~23_combout ),
	.ReadData_9(\avalonslave_0|ReadData[9]~25_combout ),
	.ReadData_15(\avalonslave_0|ReadData[15]~27_combout ),
	.ReadData_14(\avalonslave_0|ReadData[14]~29_combout ),
	.ReadData_13(\avalonslave_0|ReadData[13]~31_combout ),
	.ReadData_16(\avalonslave_0|ReadData[16]~33_combout ),
	.ReadData_20(\avalonslave_0|ReadData[20]~35_combout ),
	.ReadData_19(\avalonslave_0|ReadData[19]~37_combout ),
	.ReadData_18(\avalonslave_0|ReadData[18]~39_combout ),
	.ReadData_17(\avalonslave_0|ReadData[17]~41_combout ),
	.ReadData_23(\avalonslave_0|ReadData[23]~43_combout ),
	.ReadData_22(\avalonslave_0|ReadData[22]~45_combout ),
	.ReadData_21(\avalonslave_0|ReadData[21]~47_combout ),
	.ReadData_24(\avalonslave_0|ReadData[24]~49_combout ),
	.ReadData_31(\avalonslave_0|ReadData[31]~51_combout ),
	.ReadData_30(\avalonslave_0|ReadData[30]~53_combout ),
	.ReadData_29(\avalonslave_0|ReadData[29]~55_combout ),
	.ReadData_28(\avalonslave_0|ReadData[28]~57_combout ),
	.ReadData_27(\avalonslave_0|ReadData[27]~59_combout ),
	.ReadData_26(\avalonslave_0|ReadData[26]~61_combout ),
	.ReadData_25(\avalonslave_0|ReadData[25]~63_combout ),
	.Clk(\clk_clk~input_o ),
	.Reset(\reset_reset_n~input_o ));

nios_mcu_altera_reset_controller rst_controller(
	.r_sync_rst1(\rst_controller|r_sync_rst~q ),
	.r_early_rst1(\rst_controller|r_early_rst~q ),
	.altera_reset_synchronizer_int_chain_1(\rst_controller|alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain[1]~0_combout ),
	.clk_clk(\clk_clk~input_o ),
	.reset_reset_n(\reset_reset_n~input_o ));

nios_mcu_nios_mcu_mm_interconnect_0 mm_interconnect_0(
	.W_alu_result_12(\nios_cpu|cpu|W_alu_result[12]~q ),
	.W_alu_result_15(\nios_cpu|cpu|W_alu_result[15]~q ),
	.W_alu_result_14(\nios_cpu|cpu|W_alu_result[14]~q ),
	.W_alu_result_13(\nios_cpu|cpu|W_alu_result[13]~q ),
	.W_alu_result_11(\nios_cpu|cpu|W_alu_result[11]~q ),
	.W_alu_result_10(\nios_cpu|cpu|W_alu_result[10]~q ),
	.W_alu_result_9(\nios_cpu|cpu|W_alu_result[9]~q ),
	.W_alu_result_8(\nios_cpu|cpu|W_alu_result[8]~q ),
	.W_alu_result_7(\nios_cpu|cpu|W_alu_result[7]~q ),
	.W_alu_result_6(\nios_cpu|cpu|W_alu_result[6]~q ),
	.W_alu_result_5(\nios_cpu|cpu|W_alu_result[5]~q ),
	.W_alu_result_4(\nios_cpu|cpu|W_alu_result[4]~q ),
	.W_alu_result_3(\nios_cpu|cpu|W_alu_result[3]~q ),
	.W_alu_result_2(\nios_cpu|cpu|W_alu_result[2]~q ),
	.q_b_22(\onchip_ram|the_altsyncram|auto_generated|q_b[22] ),
	.q_b_23(\onchip_ram|the_altsyncram|auto_generated|q_b[23] ),
	.q_a_11(\onchip_ram|the_altsyncram|auto_generated|q_a[11] ),
	.q_b_11(\onchip_ram|the_altsyncram|auto_generated|q_b[11] ),
	.q_a_13(\onchip_ram|the_altsyncram|auto_generated|q_a[13] ),
	.q_b_13(\onchip_ram|the_altsyncram|auto_generated|q_b[13] ),
	.q_a_16(\onchip_ram|the_altsyncram|auto_generated|q_a[16] ),
	.q_b_16(\onchip_ram|the_altsyncram|auto_generated|q_b[16] ),
	.q_b_12(\onchip_ram|the_altsyncram|auto_generated|q_b[12] ),
	.q_a_1(\onchip_ram|the_altsyncram|auto_generated|q_a[1] ),
	.q_a_3(\onchip_ram|the_altsyncram|auto_generated|q_a[3] ),
	.q_a_5(\onchip_ram|the_altsyncram|auto_generated|q_a[5] ),
	.q_a_4(\onchip_ram|the_altsyncram|auto_generated|q_a[4] ),
	.q_b_14(\onchip_ram|the_altsyncram|auto_generated|q_b[14] ),
	.q_a_15(\onchip_ram|the_altsyncram|auto_generated|q_a[15] ),
	.q_b_15(\onchip_ram|the_altsyncram|auto_generated|q_b[15] ),
	.q_b_18(\onchip_ram|the_altsyncram|auto_generated|q_b[18] ),
	.q_b_17(\onchip_ram|the_altsyncram|auto_generated|q_b[17] ),
	.q_b_10(\onchip_ram|the_altsyncram|auto_generated|q_b[10] ),
	.q_b_9(\onchip_ram|the_altsyncram|auto_generated|q_b[9] ),
	.q_b_8(\onchip_ram|the_altsyncram|auto_generated|q_b[8] ),
	.q_a_21(\onchip_ram|the_altsyncram|auto_generated|q_a[21] ),
	.q_b_21(\onchip_ram|the_altsyncram|auto_generated|q_b[21] ),
	.q_a_19(\onchip_ram|the_altsyncram|auto_generated|q_a[19] ),
	.q_b_19(\onchip_ram|the_altsyncram|auto_generated|q_b[19] ),
	.q_a_20(\onchip_ram|the_altsyncram|auto_generated|q_a[20] ),
	.q_b_20(\onchip_ram|the_altsyncram|auto_generated|q_b[20] ),
	.readdata_0(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[0]~q ),
	.d_writedata_24(\nios_cpu|cpu|d_writedata[24]~q ),
	.d_writedata_25(\nios_cpu|cpu|d_writedata[25]~q ),
	.d_writedata_26(\nios_cpu|cpu|d_writedata[26]~q ),
	.readdata_1(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[1]~q ),
	.readdata_3(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[3]~q ),
	.readdata_2(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[2]~q ),
	.d_writedata_27(\nios_cpu|cpu|d_writedata[27]~q ),
	.d_writedata_28(\nios_cpu|cpu|d_writedata[28]~q ),
	.d_writedata_29(\nios_cpu|cpu|d_writedata[29]~q ),
	.d_writedata_30(\nios_cpu|cpu|d_writedata[30]~q ),
	.d_writedata_31(\nios_cpu|cpu|d_writedata[31]~q ),
	.d_writedata_0(\nios_cpu|cpu|d_writedata[0]~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.Equal1(\mm_interconnect_0|router|Equal1~3_combout ),
	.rst1(\jtag_uart_0|nios_mcu_jtag_uart_0_alt_jtag_atlantic|rst1~q ),
	.mem_used_1(\mm_interconnect_0|pio_0_s1_agent_rsp_fifo|mem_used[1]~q ),
	.always0(\pio_0|always0~0_combout ),
	.d_write(\nios_cpu|cpu|d_write~q ),
	.write_accepted(\mm_interconnect_0|nios_cpu_data_master_translator|write_accepted~q ),
	.wait_latency_counter_1(\mm_interconnect_0|pio_0_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|pio_0_s1_translator|wait_latency_counter[0]~q ),
	.d_writedata_1(\nios_cpu|cpu|d_writedata[1]~q ),
	.d_writedata_2(\nios_cpu|cpu|d_writedata[2]~q ),
	.d_writedata_3(\nios_cpu|cpu|d_writedata[3]~q ),
	.d_writedata_4(\nios_cpu|cpu|d_writedata[4]~q ),
	.d_writedata_5(\nios_cpu|cpu|d_writedata[5]~q ),
	.d_writedata_6(\nios_cpu|cpu|d_writedata[6]~q ),
	.d_writedata_7(\nios_cpu|cpu|d_writedata[7]~q ),
	.read_latency_shift_reg_0(\mm_interconnect_0|pio_0_s1_translator|read_latency_shift_reg[0]~q ),
	.d_read(\nios_cpu|cpu|d_read~q ),
	.read_latency_shift_reg(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg~0_combout ),
	.m0_write(\mm_interconnect_0|pio_0_s1_agent|m0_write~0_combout ),
	.mem_73_0(\mm_interconnect_0|nios_cpu_debug_mem_slave_agent_rsp_fifo|mem[0][73]~q ),
	.mem_55_0(\mm_interconnect_0|nios_cpu_debug_mem_slave_agent_rsp_fifo|mem[0][55]~q ),
	.read_latency_shift_reg_01(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_02(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg[0]~q ),
	.WideOr1(\mm_interconnect_0|rsp_mux|WideOr1~0_combout ),
	.read_latency_shift_reg_03(\mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_04(\mm_interconnect_0|onchip_ram_s2_translator|read_latency_shift_reg[0]~q ),
	.WideOr11(\mm_interconnect_0|rsp_mux|WideOr1~combout ),
	.Equal3(\mm_interconnect_0|router|Equal3~1_combout ),
	.src_channel_4(\mm_interconnect_0|router|src_channel[4]~0_combout ),
	.mem_used_11(\mm_interconnect_0|onchip_ram_s2_agent_rsp_fifo|mem_used[1]~q ),
	.saved_grant_0(\mm_interconnect_0|cmd_mux_002|saved_grant[0]~q ),
	.waitrequest(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|the_nios_mcu_nios_cpu_cpu_nios2_ocimem|waitrequest~q ),
	.mem_used_12(\mm_interconnect_0|nios_cpu_debug_mem_slave_agent_rsp_fifo|mem_used[1]~q ),
	.av_waitrequest(\jtag_uart_0|av_waitrequest~q ),
	.mem_used_13(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_agent_rsp_fifo|mem_used[1]~q ),
	.Equal2(\mm_interconnect_0|router|Equal2~0_combout ),
	.dRead(\avalonslave_0|dRead~q ),
	.always2(\mm_interconnect_0|nios_cpu_data_master_agent|always2~0_combout ),
	.m0_read(\mm_interconnect_0|avalonslave_0_avalon_slave_0_1_agent|m0_read~0_combout ),
	.m0_read1(\mm_interconnect_0|avalonslave_0_avalon_slave_0_1_agent|m0_read~1_combout ),
	.sReadCountPipelined_0(\avalonslave_0|sReadCountPipelined[0]~32_combout ),
	.nios_cpu_data_master_waitrequest(\mm_interconnect_0|nios_cpu_data_master_translator|av_waitrequest~2_combout ),
	.F_pc_10(\nios_cpu|cpu|F_pc[10]~q ),
	.F_pc_9(\nios_cpu|cpu|F_pc[9]~q ),
	.F_pc_8(\nios_cpu|cpu|F_pc[8]~q ),
	.F_pc_7(\nios_cpu|cpu|F_pc[7]~q ),
	.F_pc_6(\nios_cpu|cpu|F_pc[6]~q ),
	.F_pc_5(\nios_cpu|cpu|F_pc[5]~q ),
	.F_pc_4(\nios_cpu|cpu|F_pc[4]~q ),
	.F_pc_3(\nios_cpu|cpu|F_pc[3]~q ),
	.F_pc_2(\nios_cpu|cpu|F_pc[2]~q ),
	.F_pc_1(\nios_cpu|cpu|F_pc[1]~q ),
	.F_pc_0(\nios_cpu|cpu|F_pc[0]~q ),
	.F_pc_13(\nios_cpu|cpu|F_pc[13]~q ),
	.F_pc_12(\nios_cpu|cpu|F_pc[12]~q ),
	.F_pc_11(\nios_cpu|cpu|F_pc[11]~q ),
	.i_read(\nios_cpu|cpu|i_read~q ),
	.WideOr12(\mm_interconnect_0|cmd_mux_002|WideOr1~combout ),
	.Equal21(\avalonslave_0|Equal2~0_combout ),
	.rf_source_valid(\mm_interconnect_0|nios_cpu_debug_mem_slave_agent|rf_source_valid~1_combout ),
	.hbreak_enabled(\nios_cpu|cpu|hbreak_enabled~q ),
	.WideOr13(\mm_interconnect_0|rsp_mux|WideOr1~1_combout ),
	.av_readdata_pre_0(\mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_01(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_02(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[0]~q ),
	.src0_valid(\mm_interconnect_0|rsp_demux_002|src0_valid~0_combout ),
	.av_readdata_pre_03(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_22(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[22]~q ),
	.read_latency_shift_reg_05(\mm_interconnect_0|onchip_ram_s1_translator|read_latency_shift_reg[0]~q ),
	.src1_valid(\mm_interconnect_0|rsp_demux_002|src1_valid~0_combout ),
	.av_readdata_pre_23(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[23]~q ),
	.av_readdata_pre_24(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[24]~q ),
	.av_readdata_pre_25(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[25]~q ),
	.av_readdata_pre_26(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[26]~q ),
	.src_payload(\mm_interconnect_0|rsp_mux_001|src_payload~0_combout ),
	.av_readdata_pre_11(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[11]~q ),
	.src_payload1(\mm_interconnect_0|rsp_mux_001|src_payload~1_combout ),
	.av_readdata_pre_13(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[13]~q ),
	.src_payload2(\mm_interconnect_0|rsp_mux_001|src_payload~2_combout ),
	.av_readdata_pre_16(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[16]~q ),
	.av_readdata_pre_12(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[12]~q ),
	.src_payload3(\mm_interconnect_0|rsp_mux_001|src_payload~3_combout ),
	.av_readdata_pre_1(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[1]~q ),
	.src_payload4(\mm_interconnect_0|rsp_mux_001|src_payload~4_combout ),
	.av_readdata_pre_3(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_2(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[2]~q ),
	.src_payload5(\mm_interconnect_0|rsp_mux_001|src_payload~5_combout ),
	.av_readdata_pre_5(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[5]~q ),
	.src_payload6(\mm_interconnect_0|rsp_mux_001|src_payload~6_combout ),
	.av_readdata_pre_4(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_14(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[14]~q ),
	.src_payload7(\mm_interconnect_0|rsp_mux_001|src_payload~7_combout ),
	.av_readdata_pre_15(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_18(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[18]~q ),
	.av_readdata_pre_17(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[17]~q ),
	.av_readdata_pre_10(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_9(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_8(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_7(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_6(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[6]~q ),
	.src_payload8(\mm_interconnect_0|rsp_mux_001|src_payload~8_combout ),
	.av_readdata_pre_21(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[21]~q ),
	.src_payload9(\mm_interconnect_0|rsp_mux_001|src_payload~9_combout ),
	.av_readdata_pre_19(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[19]~q ),
	.src_payload10(\mm_interconnect_0|rsp_mux_001|src_payload~10_combout ),
	.av_readdata_pre_20(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[20]~q ),
	.src_data_46(\mm_interconnect_0|cmd_mux_002|src_data[46]~combout ),
	.av_readdata_pre_110(\mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_111(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_112(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_27(\mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_28(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_29(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_31(\mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_32(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_33(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_41(\mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_42(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_43(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_51(\mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_52(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_53(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_61(\mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_62(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_63(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_71(\mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_72(\mm_interconnect_0|jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_73(\mm_interconnect_0|pio_0_s1_translator|av_readdata_pre[7]~q ),
	.b_full(\jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.src_data_8(\mm_interconnect_0|rsp_mux|src_data[8]~1_combout ),
	.ReadData_0(\avalonslave_0|ReadData[0]~1_combout ),
	.read_0(\jtag_uart_0|read_0~q ),
	.av_readdata_0(\jtag_uart_0|av_readdata[0]~0_combout ),
	.d_byteenable_0(\nios_cpu|cpu|d_byteenable[0]~q ),
	.readdata_01(\pio_0|readdata[0]~combout ),
	.av_readdata_9(\jtag_uart_0|av_readdata[9]~combout ),
	.av_readdata_8(\jtag_uart_0|av_readdata[8]~1_combout ),
	.readdata_22(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[22]~q ),
	.d_writedata_22(\nios_cpu|cpu|d_writedata[22]~q ),
	.d_byteenable_2(\nios_cpu|cpu|d_byteenable[2]~q ),
	.readdata_23(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[23]~q ),
	.d_writedata_23(\nios_cpu|cpu|d_writedata[23]~q ),
	.readdata_24(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[24]~q ),
	.d_byteenable_3(\nios_cpu|cpu|d_byteenable[3]~q ),
	.readdata_25(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[25]~q ),
	.readdata_26(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[26]~q ),
	.d_writedata_11(\nios_cpu|cpu|d_writedata[11]~q ),
	.d_byteenable_1(\nios_cpu|cpu|d_byteenable[1]~q ),
	.readdata_11(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[11]~q ),
	.d_writedata_13(\nios_cpu|cpu|d_writedata[13]~q ),
	.readdata_13(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[13]~q ),
	.d_writedata_16(\nios_cpu|cpu|d_writedata[16]~q ),
	.readdata_16(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[16]~q ),
	.readdata_12(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[12]~q ),
	.d_writedata_12(\nios_cpu|cpu|d_writedata[12]~q ),
	.readdata_5(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[5]~q ),
	.readdata_4(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[4]~q ),
	.d_writedata_14(\nios_cpu|cpu|d_writedata[14]~q ),
	.readdata_14(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[14]~q ),
	.d_writedata_15(\nios_cpu|cpu|d_writedata[15]~q ),
	.readdata_15(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[15]~q ),
	.d_writedata_18(\nios_cpu|cpu|d_writedata[18]~q ),
	.readdata_18(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[18]~q ),
	.src_data_12(\mm_interconnect_0|rsp_mux|src_data[12]~3_combout ),
	.av_readdata_pre_271(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[27]~q ),
	.av_readdata_pre_281(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[28]~q ),
	.av_readdata_pre_291(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[29]~q ),
	.av_readdata_pre_30(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[30]~q ),
	.av_readdata_pre_311(\mm_interconnect_0|nios_cpu_debug_mem_slave_translator|av_readdata_pre[31]~q ),
	.d_writedata_17(\nios_cpu|cpu|d_writedata[17]~q ),
	.readdata_17(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[17]~q ),
	.src_data_11(\mm_interconnect_0|rsp_mux|src_data[11]~combout ),
	.src_data_10(\mm_interconnect_0|rsp_mux|src_data[10]~6_combout ),
	.src_data_9(\mm_interconnect_0|rsp_mux|src_data[9]~8_combout ),
	.readdata_10(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[10]~q ),
	.d_writedata_10(\nios_cpu|cpu|d_writedata[10]~q ),
	.readdata_9(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[9]~q ),
	.d_writedata_9(\nios_cpu|cpu|d_writedata[9]~q ),
	.readdata_8(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[8]~q ),
	.d_writedata_8(\nios_cpu|cpu|d_writedata[8]~q ),
	.readdata_7(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[7]~q ),
	.readdata_6(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[6]~q ),
	.d_writedata_21(\nios_cpu|cpu|d_writedata[21]~q ),
	.readdata_21(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[21]~q ),
	.src_data_15(\mm_interconnect_0|rsp_mux|src_data[15]~10_combout ),
	.d_writedata_19(\nios_cpu|cpu|d_writedata[19]~q ),
	.readdata_19(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[19]~q ),
	.d_writedata_20(\nios_cpu|cpu|d_writedata[20]~q ),
	.readdata_20(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[20]~q ),
	.src_data_14(\mm_interconnect_0|rsp_mux|src_data[14]~12_combout ),
	.src_data_13(\mm_interconnect_0|rsp_mux|src_data[13]~14_combout ),
	.ReadData_1(\avalonslave_0|ReadData[1]~3_combout ),
	.av_readdata_1(\jtag_uart_0|av_readdata[1]~2_combout ),
	.readdata_110(\pio_0|readdata[1]~combout ),
	.ReadData_2(\avalonslave_0|ReadData[2]~5_combout ),
	.av_readdata_2(\jtag_uart_0|av_readdata[2]~3_combout ),
	.readdata_27(\pio_0|readdata[2]~combout ),
	.ReadData_3(\avalonslave_0|ReadData[3]~7_combout ),
	.av_readdata_3(\jtag_uart_0|av_readdata[3]~4_combout ),
	.readdata_31(\pio_0|readdata[3]~combout ),
	.ReadData_4(\avalonslave_0|ReadData[4]~9_combout ),
	.av_readdata_4(\jtag_uart_0|av_readdata[4]~5_combout ),
	.readdata_41(\pio_0|readdata[4]~combout ),
	.ReadData_5(\avalonslave_0|ReadData[5]~11_combout ),
	.av_readdata_5(\jtag_uart_0|av_readdata[5]~6_combout ),
	.readdata_51(\pio_0|readdata[5]~combout ),
	.ReadData_6(\avalonslave_0|ReadData[6]~13_combout ),
	.av_readdata_6(\jtag_uart_0|av_readdata[6]~7_combout ),
	.readdata_61(\pio_0|readdata[6]~combout ),
	.ReadData_7(\avalonslave_0|ReadData[7]~15_combout ),
	.av_readdata_7(\jtag_uart_0|av_readdata[7]~8_combout ),
	.readdata_71(\pio_0|readdata[7]~combout ),
	.b_non_empty(\jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.counter_reg_bit_5(\jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.counter_reg_bit_4(\jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.counter_reg_bit_2(\jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.src_payload11(\mm_interconnect_0|cmd_mux_002|src_payload~0_combout ),
	.src_payload12(\mm_interconnect_0|cmd_mux_002|src_payload~1_combout ),
	.src_data_38(\mm_interconnect_0|cmd_mux_002|src_data[38]~combout ),
	.src_data_39(\mm_interconnect_0|cmd_mux_002|src_data[39]~combout ),
	.src_data_40(\mm_interconnect_0|cmd_mux_002|src_data[40]~combout ),
	.src_data_41(\mm_interconnect_0|cmd_mux_002|src_data[41]~combout ),
	.src_data_42(\mm_interconnect_0|cmd_mux_002|src_data[42]~combout ),
	.src_data_43(\mm_interconnect_0|cmd_mux_002|src_data[43]~combout ),
	.src_data_44(\mm_interconnect_0|cmd_mux_002|src_data[44]~combout ),
	.src_data_45(\mm_interconnect_0|cmd_mux_002|src_data[45]~combout ),
	.src_data_32(\mm_interconnect_0|cmd_mux_002|src_data[32]~combout ),
	.ReadData_8(\avalonslave_0|ReadData[8]~17_combout ),
	.src_data_16(\mm_interconnect_0|rsp_mux|src_data[16]~16_combout ),
	.counter_reg_bit_31(\jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.counter_reg_bit_01(\jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.counter_reg_bit_21(\jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.counter_reg_bit_11(\jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.b_full1(\jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.counter_reg_bit_51(\jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.counter_reg_bit_41(\jtag_uart_0|the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.ReadData_12(\avalonslave_0|ReadData[12]~19_combout ),
	.src_data_20(\mm_interconnect_0|rsp_mux|src_data[20]~18_combout ),
	.readdata_271(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[27]~q ),
	.readdata_28(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[28]~q ),
	.readdata_29(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[29]~q ),
	.readdata_30(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[30]~q ),
	.readdata_311(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|readdata[31]~q ),
	.ReadData_11(\avalonslave_0|ReadData[11]~21_combout ),
	.src_data_19(\mm_interconnect_0|rsp_mux|src_data[19]~20_combout ),
	.ReadData_10(\avalonslave_0|ReadData[10]~23_combout ),
	.ac(\jtag_uart_0|ac~q ),
	.src_data_18(\mm_interconnect_0|rsp_mux|src_data[18]~22_combout ),
	.ReadData_9(\avalonslave_0|ReadData[9]~25_combout ),
	.src_data_17(\mm_interconnect_0|rsp_mux|src_data[17]~24_combout ),
	.ReadData_15(\avalonslave_0|ReadData[15]~27_combout ),
	.rvalid(\jtag_uart_0|rvalid~q ),
	.src_data_23(\mm_interconnect_0|rsp_mux|src_data[23]~combout ),
	.ReadData_14(\avalonslave_0|ReadData[14]~29_combout ),
	.woverflow(\jtag_uart_0|woverflow~q ),
	.src_data_22(\mm_interconnect_0|rsp_mux|src_data[22]~27_combout ),
	.ReadData_13(\avalonslave_0|ReadData[13]~31_combout ),
	.src_data_21(\mm_interconnect_0|rsp_mux|src_data[21]~29_combout ),
	.src_payload13(\mm_interconnect_0|cmd_mux_002|src_payload~2_combout ),
	.ReadData_16(\avalonslave_0|ReadData[16]~33_combout ),
	.av_readdata_pre_241(\mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[24]~q ),
	.av_readdata_pre_312(\mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[31]~q ),
	.av_readdata_pre_301(\mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[30]~q ),
	.av_readdata_pre_292(\mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[29]~q ),
	.av_readdata_pre_282(\mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[28]~q ),
	.av_readdata_pre_272(\mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[27]~q ),
	.av_readdata_pre_261(\mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[26]~q ),
	.av_readdata_pre_251(\mm_interconnect_0|avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[25]~q ),
	.src_payload14(\mm_interconnect_0|cmd_mux_002|src_payload~3_combout ),
	.ReadData_20(\avalonslave_0|ReadData[20]~35_combout ),
	.ReadData_19(\avalonslave_0|ReadData[19]~37_combout ),
	.ReadData_18(\avalonslave_0|ReadData[18]~39_combout ),
	.ReadData_17(\avalonslave_0|ReadData[17]~41_combout ),
	.ReadData_23(\avalonslave_0|ReadData[23]~43_combout ),
	.ReadData_22(\avalonslave_0|ReadData[22]~45_combout ),
	.ReadData_21(\avalonslave_0|ReadData[21]~47_combout ),
	.src_payload15(\mm_interconnect_0|cmd_mux_002|src_payload~4_combout ),
	.ReadData_24(\avalonslave_0|ReadData[24]~49_combout ),
	.ReadData_31(\avalonslave_0|ReadData[31]~51_combout ),
	.ReadData_30(\avalonslave_0|ReadData[30]~53_combout ),
	.ReadData_29(\avalonslave_0|ReadData[29]~55_combout ),
	.ReadData_28(\avalonslave_0|ReadData[28]~57_combout ),
	.ReadData_27(\avalonslave_0|ReadData[27]~59_combout ),
	.ReadData_26(\avalonslave_0|ReadData[26]~61_combout ),
	.ReadData_25(\avalonslave_0|ReadData[25]~63_combout ),
	.src_payload16(\mm_interconnect_0|cmd_mux_002|src_payload~5_combout ),
	.src_data_34(\mm_interconnect_0|cmd_mux_002|src_data[34]~combout ),
	.src_payload17(\mm_interconnect_0|cmd_mux_002|src_payload~6_combout ),
	.src_payload18(\mm_interconnect_0|cmd_mux_002|src_payload~7_combout ),
	.src_data_35(\mm_interconnect_0|cmd_mux_002|src_data[35]~combout ),
	.src_payload19(\mm_interconnect_0|cmd_mux_002|src_payload~8_combout ),
	.src_payload20(\mm_interconnect_0|cmd_mux_002|src_payload~9_combout ),
	.src_payload21(\mm_interconnect_0|cmd_mux_002|src_payload~10_combout ),
	.src_data_33(\mm_interconnect_0|cmd_mux_002|src_data[33]~combout ),
	.src_payload22(\mm_interconnect_0|cmd_mux_002|src_payload~11_combout ),
	.src_payload23(\mm_interconnect_0|cmd_mux_002|src_payload~12_combout ),
	.src_payload24(\mm_interconnect_0|cmd_mux_002|src_payload~13_combout ),
	.src_payload25(\mm_interconnect_0|cmd_mux_002|src_payload~14_combout ),
	.src_payload26(\mm_interconnect_0|cmd_mux_002|src_payload~15_combout ),
	.src_payload27(\mm_interconnect_0|cmd_mux_002|src_payload~16_combout ),
	.src_payload28(\mm_interconnect_0|cmd_mux_002|src_payload~17_combout ),
	.src_payload29(\mm_interconnect_0|cmd_mux_002|src_payload~18_combout ),
	.src_payload30(\mm_interconnect_0|cmd_mux_002|src_payload~19_combout ),
	.src_payload31(\mm_interconnect_0|cmd_mux_002|src_payload~20_combout ),
	.src_payload32(\mm_interconnect_0|cmd_mux_002|src_payload~21_combout ),
	.src_payload33(\mm_interconnect_0|cmd_mux_002|src_payload~22_combout ),
	.src_payload34(\mm_interconnect_0|cmd_mux_002|src_payload~23_combout ),
	.src_payload35(\mm_interconnect_0|cmd_mux_002|src_payload~24_combout ),
	.src_payload36(\mm_interconnect_0|cmd_mux_002|src_payload~25_combout ),
	.src_payload37(\mm_interconnect_0|cmd_mux_002|src_payload~26_combout ),
	.src_payload38(\mm_interconnect_0|cmd_mux_002|src_payload~27_combout ),
	.src_payload39(\mm_interconnect_0|cmd_mux_002|src_payload~28_combout ),
	.src_payload40(\mm_interconnect_0|cmd_mux_002|src_payload~29_combout ),
	.src_payload41(\mm_interconnect_0|cmd_mux_002|src_payload~30_combout ),
	.src_payload42(\mm_interconnect_0|cmd_mux_002|src_payload~31_combout ),
	.src_payload43(\mm_interconnect_0|cmd_mux_002|src_payload~32_combout ),
	.clk_clk(\clk_clk~input_o ));

nios_mcu_nios_mcu_pio_0 pio_0(
	.W_alu_result_4(\nios_cpu|cpu|W_alu_result[4]~q ),
	.W_alu_result_3(\nios_cpu|cpu|W_alu_result[3]~q ),
	.W_alu_result_2(\nios_cpu|cpu|W_alu_result[2]~q ),
	.data_out_0(\pio_0|data_out[0]~q ),
	.data_out_1(\pio_0|data_out[1]~q ),
	.data_out_2(\pio_0|data_out[2]~q ),
	.data_out_3(\pio_0|data_out[3]~q ),
	.data_out_4(\pio_0|data_out[4]~q ),
	.data_out_5(\pio_0|data_out[5]~q ),
	.data_out_6(\pio_0|data_out[6]~q ),
	.data_out_7(\pio_0|data_out[7]~q ),
	.writedata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\nios_cpu|cpu|d_writedata[7]~q ,\nios_cpu|cpu|d_writedata[6]~q ,\nios_cpu|cpu|d_writedata[5]~q ,\nios_cpu|cpu|d_writedata[4]~q ,\nios_cpu|cpu|d_writedata[3]~q ,
\nios_cpu|cpu|d_writedata[2]~q ,\nios_cpu|cpu|d_writedata[1]~q ,\nios_cpu|cpu|d_writedata[0]~q }),
	.reset_n(\rst_controller|r_sync_rst~q ),
	.Equal1(\mm_interconnect_0|router|Equal1~3_combout ),
	.rst1(\jtag_uart_0|nios_mcu_jtag_uart_0_alt_jtag_atlantic|rst1~q ),
	.mem_used_1(\mm_interconnect_0|pio_0_s1_agent_rsp_fifo|mem_used[1]~q ),
	.always0(\pio_0|always0~0_combout ),
	.d_write(\nios_cpu|cpu|d_write~q ),
	.write_accepted(\mm_interconnect_0|nios_cpu_data_master_translator|write_accepted~q ),
	.wait_latency_counter_1(\mm_interconnect_0|pio_0_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|pio_0_s1_translator|wait_latency_counter[0]~q ),
	.readdata_0(\pio_0|readdata[0]~combout ),
	.readdata_1(\pio_0|readdata[1]~combout ),
	.readdata_2(\pio_0|readdata[2]~combout ),
	.readdata_3(\pio_0|readdata[3]~combout ),
	.readdata_4(\pio_0|readdata[4]~combout ),
	.readdata_5(\pio_0|readdata[5]~combout ),
	.readdata_6(\pio_0|readdata[6]~combout ),
	.readdata_7(\pio_0|readdata[7]~combout ),
	.clk(\clk_clk~input_o ));

nios_mcu_nios_mcu_onchip_ram onchip_ram(
	.W_alu_result_12(\nios_cpu|cpu|W_alu_result[12]~q ),
	.W_alu_result_14(\nios_cpu|cpu|W_alu_result[14]~q ),
	.W_alu_result_13(\nios_cpu|cpu|W_alu_result[13]~q ),
	.W_alu_result_11(\nios_cpu|cpu|W_alu_result[11]~q ),
	.W_alu_result_10(\nios_cpu|cpu|W_alu_result[10]~q ),
	.W_alu_result_9(\nios_cpu|cpu|W_alu_result[9]~q ),
	.W_alu_result_8(\nios_cpu|cpu|W_alu_result[8]~q ),
	.W_alu_result_7(\nios_cpu|cpu|W_alu_result[7]~q ),
	.W_alu_result_6(\nios_cpu|cpu|W_alu_result[6]~q ),
	.W_alu_result_5(\nios_cpu|cpu|W_alu_result[5]~q ),
	.W_alu_result_4(\nios_cpu|cpu|W_alu_result[4]~q ),
	.W_alu_result_3(\nios_cpu|cpu|W_alu_result[3]~q ),
	.W_alu_result_2(\nios_cpu|cpu|W_alu_result[2]~q ),
	.q_a_0(\onchip_ram|the_altsyncram|auto_generated|q_a[0] ),
	.q_b_0(\onchip_ram|the_altsyncram|auto_generated|q_b[0] ),
	.q_a_22(\onchip_ram|the_altsyncram|auto_generated|q_a[22] ),
	.q_b_22(\onchip_ram|the_altsyncram|auto_generated|q_b[22] ),
	.q_a_23(\onchip_ram|the_altsyncram|auto_generated|q_a[23] ),
	.q_b_23(\onchip_ram|the_altsyncram|auto_generated|q_b[23] ),
	.q_a_24(\onchip_ram|the_altsyncram|auto_generated|q_a[24] ),
	.q_b_24(\onchip_ram|the_altsyncram|auto_generated|q_b[24] ),
	.q_a_25(\onchip_ram|the_altsyncram|auto_generated|q_a[25] ),
	.q_b_25(\onchip_ram|the_altsyncram|auto_generated|q_b[25] ),
	.q_a_26(\onchip_ram|the_altsyncram|auto_generated|q_a[26] ),
	.q_b_26(\onchip_ram|the_altsyncram|auto_generated|q_b[26] ),
	.q_a_11(\onchip_ram|the_altsyncram|auto_generated|q_a[11] ),
	.q_b_11(\onchip_ram|the_altsyncram|auto_generated|q_b[11] ),
	.q_a_13(\onchip_ram|the_altsyncram|auto_generated|q_a[13] ),
	.q_b_13(\onchip_ram|the_altsyncram|auto_generated|q_b[13] ),
	.q_a_16(\onchip_ram|the_altsyncram|auto_generated|q_a[16] ),
	.q_b_16(\onchip_ram|the_altsyncram|auto_generated|q_b[16] ),
	.q_a_12(\onchip_ram|the_altsyncram|auto_generated|q_a[12] ),
	.q_b_12(\onchip_ram|the_altsyncram|auto_generated|q_b[12] ),
	.q_a_1(\onchip_ram|the_altsyncram|auto_generated|q_a[1] ),
	.q_b_1(\onchip_ram|the_altsyncram|auto_generated|q_b[1] ),
	.q_a_3(\onchip_ram|the_altsyncram|auto_generated|q_a[3] ),
	.q_b_3(\onchip_ram|the_altsyncram|auto_generated|q_b[3] ),
	.q_a_2(\onchip_ram|the_altsyncram|auto_generated|q_a[2] ),
	.q_b_2(\onchip_ram|the_altsyncram|auto_generated|q_b[2] ),
	.q_a_5(\onchip_ram|the_altsyncram|auto_generated|q_a[5] ),
	.q_b_5(\onchip_ram|the_altsyncram|auto_generated|q_b[5] ),
	.q_a_4(\onchip_ram|the_altsyncram|auto_generated|q_a[4] ),
	.q_b_4(\onchip_ram|the_altsyncram|auto_generated|q_b[4] ),
	.q_a_14(\onchip_ram|the_altsyncram|auto_generated|q_a[14] ),
	.q_b_14(\onchip_ram|the_altsyncram|auto_generated|q_b[14] ),
	.q_a_15(\onchip_ram|the_altsyncram|auto_generated|q_a[15] ),
	.q_b_15(\onchip_ram|the_altsyncram|auto_generated|q_b[15] ),
	.q_a_18(\onchip_ram|the_altsyncram|auto_generated|q_a[18] ),
	.q_b_18(\onchip_ram|the_altsyncram|auto_generated|q_b[18] ),
	.q_a_17(\onchip_ram|the_altsyncram|auto_generated|q_a[17] ),
	.q_b_17(\onchip_ram|the_altsyncram|auto_generated|q_b[17] ),
	.q_a_10(\onchip_ram|the_altsyncram|auto_generated|q_a[10] ),
	.q_b_10(\onchip_ram|the_altsyncram|auto_generated|q_b[10] ),
	.q_a_9(\onchip_ram|the_altsyncram|auto_generated|q_a[9] ),
	.q_b_9(\onchip_ram|the_altsyncram|auto_generated|q_b[9] ),
	.q_a_8(\onchip_ram|the_altsyncram|auto_generated|q_a[8] ),
	.q_b_8(\onchip_ram|the_altsyncram|auto_generated|q_b[8] ),
	.q_a_7(\onchip_ram|the_altsyncram|auto_generated|q_a[7] ),
	.q_b_7(\onchip_ram|the_altsyncram|auto_generated|q_b[7] ),
	.q_a_6(\onchip_ram|the_altsyncram|auto_generated|q_a[6] ),
	.q_b_6(\onchip_ram|the_altsyncram|auto_generated|q_b[6] ),
	.q_a_21(\onchip_ram|the_altsyncram|auto_generated|q_a[21] ),
	.q_b_21(\onchip_ram|the_altsyncram|auto_generated|q_b[21] ),
	.q_a_19(\onchip_ram|the_altsyncram|auto_generated|q_a[19] ),
	.q_b_19(\onchip_ram|the_altsyncram|auto_generated|q_b[19] ),
	.q_a_20(\onchip_ram|the_altsyncram|auto_generated|q_a[20] ),
	.q_b_20(\onchip_ram|the_altsyncram|auto_generated|q_b[20] ),
	.d_writedata_24(\nios_cpu|cpu|d_writedata[24]~q ),
	.d_writedata_25(\nios_cpu|cpu|d_writedata[25]~q ),
	.d_writedata_26(\nios_cpu|cpu|d_writedata[26]~q ),
	.q_a_27(\onchip_ram|the_altsyncram|auto_generated|q_a[27] ),
	.q_b_27(\onchip_ram|the_altsyncram|auto_generated|q_b[27] ),
	.q_a_28(\onchip_ram|the_altsyncram|auto_generated|q_a[28] ),
	.q_b_28(\onchip_ram|the_altsyncram|auto_generated|q_b[28] ),
	.q_a_29(\onchip_ram|the_altsyncram|auto_generated|q_a[29] ),
	.q_b_29(\onchip_ram|the_altsyncram|auto_generated|q_b[29] ),
	.q_a_30(\onchip_ram|the_altsyncram|auto_generated|q_a[30] ),
	.q_b_30(\onchip_ram|the_altsyncram|auto_generated|q_b[30] ),
	.q_a_31(\onchip_ram|the_altsyncram|auto_generated|q_a[31] ),
	.q_b_31(\onchip_ram|the_altsyncram|auto_generated|q_b[31] ),
	.d_writedata_27(\nios_cpu|cpu|d_writedata[27]~q ),
	.d_writedata_28(\nios_cpu|cpu|d_writedata[28]~q ),
	.d_writedata_29(\nios_cpu|cpu|d_writedata[29]~q ),
	.d_writedata_30(\nios_cpu|cpu|d_writedata[30]~q ),
	.d_writedata_31(\nios_cpu|cpu|d_writedata[31]~q ),
	.d_writedata_0(\nios_cpu|cpu|d_writedata[0]~q ),
	.rst1(\jtag_uart_0|nios_mcu_jtag_uart_0_alt_jtag_atlantic|rst1~q ),
	.d_writedata_1(\nios_cpu|cpu|d_writedata[1]~q ),
	.d_writedata_2(\nios_cpu|cpu|d_writedata[2]~q ),
	.d_writedata_3(\nios_cpu|cpu|d_writedata[3]~q ),
	.d_writedata_4(\nios_cpu|cpu|d_writedata[4]~q ),
	.d_writedata_5(\nios_cpu|cpu|d_writedata[5]~q ),
	.d_writedata_6(\nios_cpu|cpu|d_writedata[6]~q ),
	.d_writedata_7(\nios_cpu|cpu|d_writedata[7]~q ),
	.m0_write(\mm_interconnect_0|pio_0_s1_agent|m0_write~0_combout ),
	.src_channel_4(\mm_interconnect_0|router|src_channel[4]~0_combout ),
	.mem_used_1(\mm_interconnect_0|onchip_ram_s2_agent_rsp_fifo|mem_used[1]~q ),
	.F_pc_10(\nios_cpu|cpu|F_pc[10]~q ),
	.F_pc_9(\nios_cpu|cpu|F_pc[9]~q ),
	.F_pc_8(\nios_cpu|cpu|F_pc[8]~q ),
	.F_pc_7(\nios_cpu|cpu|F_pc[7]~q ),
	.F_pc_6(\nios_cpu|cpu|F_pc[6]~q ),
	.F_pc_5(\nios_cpu|cpu|F_pc[5]~q ),
	.F_pc_4(\nios_cpu|cpu|F_pc[4]~q ),
	.F_pc_3(\nios_cpu|cpu|F_pc[3]~q ),
	.F_pc_2(\nios_cpu|cpu|F_pc[2]~q ),
	.F_pc_1(\nios_cpu|cpu|F_pc[1]~q ),
	.F_pc_0(\nios_cpu|cpu|F_pc[0]~q ),
	.F_pc_12(\nios_cpu|cpu|F_pc[12]~q ),
	.F_pc_11(\nios_cpu|cpu|F_pc[11]~q ),
	.r_early_rst(\rst_controller|r_early_rst~q ),
	.d_byteenable_0(\nios_cpu|cpu|d_byteenable[0]~q ),
	.d_writedata_22(\nios_cpu|cpu|d_writedata[22]~q ),
	.d_byteenable_2(\nios_cpu|cpu|d_byteenable[2]~q ),
	.d_writedata_23(\nios_cpu|cpu|d_writedata[23]~q ),
	.d_byteenable_3(\nios_cpu|cpu|d_byteenable[3]~q ),
	.d_writedata_11(\nios_cpu|cpu|d_writedata[11]~q ),
	.d_byteenable_1(\nios_cpu|cpu|d_byteenable[1]~q ),
	.d_writedata_13(\nios_cpu|cpu|d_writedata[13]~q ),
	.d_writedata_16(\nios_cpu|cpu|d_writedata[16]~q ),
	.d_writedata_12(\nios_cpu|cpu|d_writedata[12]~q ),
	.d_writedata_14(\nios_cpu|cpu|d_writedata[14]~q ),
	.d_writedata_15(\nios_cpu|cpu|d_writedata[15]~q ),
	.d_writedata_18(\nios_cpu|cpu|d_writedata[18]~q ),
	.d_writedata_17(\nios_cpu|cpu|d_writedata[17]~q ),
	.d_writedata_10(\nios_cpu|cpu|d_writedata[10]~q ),
	.d_writedata_9(\nios_cpu|cpu|d_writedata[9]~q ),
	.d_writedata_8(\nios_cpu|cpu|d_writedata[8]~q ),
	.d_writedata_21(\nios_cpu|cpu|d_writedata[21]~q ),
	.d_writedata_19(\nios_cpu|cpu|d_writedata[19]~q ),
	.d_writedata_20(\nios_cpu|cpu|d_writedata[20]~q ),
	.GND_port(\~GND~combout ),
	.clk_clk(\clk_clk~input_o ));

cycloneive_lcell_comb \~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\~GND~combout ),
	.cout());
defparam \~GND .lut_mask = 16'h0000;
defparam \~GND .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~4_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~6_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~4_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~7_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~9_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~10_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~9_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 (
	.dataa(gnd),
	.datab(\altera_internal_jtag~TMSUTAP ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .lut_mask = 16'h3FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.datab(\altera_internal_jtag~TDIUTAP ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .lut_mask = 16'hFFF7;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~4 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(\altera_internal_jtag~TDIUTAP ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~5 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~5_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~6 .lut_mask = 16'hFFF7;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~6 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~6_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~7_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~7 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0 .lut_mask = 16'hEEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~8 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~8_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~1_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~9 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~9 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~8_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~7_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~10 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~1 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~6 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~1_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~7 .lut_mask = 16'hFAFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~8 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~8 .sum_lutc_input = "datac";

assign \clk_clk~input_o  = clk_clk;

assign \reset_reset_n~input_o  = reset_reset_n;

assign leds_export[0] = \pio_0|data_out[0]~q ;

assign leds_export[1] = \pio_0|data_out[1]~q ;

assign leds_export[2] = \pio_0|data_out[2]~q ;

assign leds_export[3] = \pio_0|data_out[3]~q ;

assign leds_export[4] = \pio_0|data_out[4]~q ;

assign leds_export[5] = \pio_0|data_out[5]~q ;

assign leds_export[6] = \pio_0|data_out[6]~q ;

assign leds_export[7] = \pio_0|data_out[7]~q ;

assign altera_reserved_tdo = \altera_internal_jtag~TDO ;

assign \altera_reserved_tms~input_o  = altera_reserved_tms;

assign \altera_reserved_tck~input_o  = altera_reserved_tck;

assign \altera_reserved_tdi~input_o  = altera_reserved_tdi;

cycloneive_jtag altera_internal_jtag(
	.tms(\altera_reserved_tms~input_o ),
	.tck(\altera_reserved_tck~input_o ),
	.tdi(\altera_reserved_tdi~input_o ),
	.tdoutap(gnd),
	.tdouser(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.tdo(\altera_internal_jtag~TDO ),
	.tmsutap(\altera_internal_jtag~TMSUTAP ),
	.tckutap(\altera_internal_jtag~TCKUTAP ),
	.tdiutap(\altera_internal_jtag~TDIUTAP ),
	.shiftuser(),
	.clkdruser(),
	.updateuser(),
	.runidleuser(),
	.usr1user());

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\altera_internal_jtag~TMSUTAP ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .lut_mask = 16'h0FF0;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 (
	.dataa(gnd),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .lut_mask = 16'hC33C;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .lut_mask = 16'hFF7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\altera_internal_jtag~TMSUTAP ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .lut_mask = 16'h7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 .lut_mask = 16'hEEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\rst_controller|alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain[1]~0_combout ),
	.datac(\rst_controller|alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain[1]~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~6 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 (
	.dataa(\altera_internal_jtag~TDIUTAP ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~6_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~7 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~7_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~14 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~14_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~14 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~9 (
	.dataa(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_tck|ir_out[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~9 .lut_mask = 16'hFAFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~9 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~9_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~16_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~7 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~7 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~7_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~10 .lut_mask = 16'hFFB8;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~16 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~10_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~16_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~16 .lut_mask = 16'hFFAC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~16 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~14_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~16_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~15 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~15_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~15 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~15 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~15_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~16_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~13 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~13 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~13_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~16_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0 (
	.dataa(gnd),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0 .lut_mask = 16'h3FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~8 .lut_mask = 16'hF7FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~3 .lut_mask = 16'h8B8B;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~8_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~3_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~4 .lut_mask = 16'hB8FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~4 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~4_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~14_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~5 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~5 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~1 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~1_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 .lut_mask = 16'hFAFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~3 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~3_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~4 .lut_mask = 16'hFFAC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~5 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~4_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~5_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~6 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~6 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~6_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~11_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~11 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~12 (
	.dataa(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_tck|ir_out[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~11_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~12_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~12 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~12 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~12_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~16_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~6 .lut_mask = 16'hFAFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~6 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~6_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~4 .lut_mask = 16'hEEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~4_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 (
	.dataa(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(\jtag_uart_0|nios_mcu_jtag_uart_0_alt_jtag_atlantic|adapted_tdo~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 .lut_mask = 16'hFAFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~9_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~10 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~9 .lut_mask = 16'h55AA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~12 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~10 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~12_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~13 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~12 .lut_mask = 16'h5A5F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~11_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~11 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~11 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~20_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~11_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~14 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~13 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~14_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~15 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~14 .lut_mask = 16'h5AAF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~14 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~20_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~11_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~16 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~15 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~16_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~17 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~16 .lut_mask = 16'h5A5F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~16 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~20_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~11_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~18 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~17 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~18_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~18 .lut_mask = 16'h5A5A;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~18 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~20_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~11_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~20 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~16_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~20_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~20 .lut_mask = 16'hFFF7;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~20 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~20_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~11_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~16 (
	.dataa(gnd),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~16_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~16 .lut_mask = 16'h3FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~17 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~17_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~17 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~18 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~16_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~17_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~18_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~18 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~19 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~19_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~19 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~20 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~19_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~20_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~20 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~18_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~20_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~25 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~25_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~25 .lut_mask = 16'h6996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~26 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~25_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~26_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~26 .lut_mask = 16'hF7FD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~26 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~26_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~20_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~23 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~23_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~23 .lut_mask = 16'h6996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~24 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~23_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~24_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~24 .lut_mask = 16'hCF5F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~24 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~24_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~20_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~21 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~21_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~21 .lut_mask = 16'hD77D;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~22 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~21_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~22_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~22 .lut_mask = 16'h9F6F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~22 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~22_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~20_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .lut_mask = 16'h0FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena (
	.dataa(gnd),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena .lut_mask = 16'hFFFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3_combout ),
	.asdata(\altera_internal_jtag~TDIUTAP ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~12 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11 .lut_mask = 16'h55AA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~17 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~17_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~17 .lut_mask = 16'h5A5F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~17 .sum_lutc_input = "cin";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20 .lut_mask = 16'h5A5A;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20 .sum_lutc_input = "cin";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~23 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~23_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~23 .lut_mask = 16'hFFFB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~23 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~19 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~19_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~19 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~22 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~19_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~22_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~22 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~22 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~12 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~14 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13 .lut_mask = 16'h5A5F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~15 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~14 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~15_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~15 .lut_mask = 16'h5AAF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~15 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .lut_mask = 16'h7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datab(gnd),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~13 .lut_mask = 16'hAFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~14 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~13_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~14_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~14 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~16 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~16_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~16 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~17 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~16_combout ),
	.datab(\altera_internal_jtag~TDIUTAP ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~17_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~17 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~19 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~19_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~19 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~19 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~19_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~15 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~14_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~15_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~15 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~15 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~19_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~19_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~18 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~18_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~18 .lut_mask = 16'hFFF7;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 .lut_mask = 16'h6996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~18_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 .lut_mask = 16'hEFEF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~19_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .lut_mask = 16'hFFBE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .lut_mask = 16'hFFDF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 (
	.dataa(\jtag_uart_0|nios_mcu_jtag_uart_0_alt_jtag_atlantic|adapted_tdo~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .lut_mask = 16'hACFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ),
	.datab(\nios_cpu|cpu|the_nios_mcu_nios_cpu_cpu_nios2_oci|the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 (
	.dataa(\altera_internal_jtag~TDIUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datab(gnd),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~8 .lut_mask = 16'hAFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~8_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~9 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~9_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~10 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~10 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo (
	.clk(!\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .power_up = "low";

cycloneive_lcell_comb \auto_hub|~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|~GND~combout ),
	.cout());
defparam \auto_hub|~GND .lut_mask = 16'h0000;
defparam \auto_hub|~GND .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .sum_lutc_input = "datac";

endmodule

module nios_mcu_altera_reset_controller (
	r_sync_rst1,
	r_early_rst1,
	altera_reset_synchronizer_int_chain_1,
	clk_clk,
	reset_reset_n)/* synthesis synthesis_greybox=1 */;
output 	r_sync_rst1;
output 	r_early_rst1;
output 	altera_reset_synchronizer_int_chain_1;
input 	clk_clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;
wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[2]~q ;
wire \altera_reset_synchronizer_int_chain[3]~q ;
wire \altera_reset_synchronizer_int_chain[4]~0_combout ;
wire \altera_reset_synchronizer_int_chain[4]~q ;
wire \r_sync_rst_chain[3]~q ;
wire \r_sync_rst_chain~1_combout ;
wire \r_sync_rst_chain[2]~q ;
wire \r_sync_rst_chain~0_combout ;
wire \r_sync_rst_chain[1]~q ;
wire \WideOr0~0_combout ;
wire \always2~0_combout ;


nios_mcu_altera_reset_synchronizer alt_rst_req_sync_uq1(
	.altera_reset_synchronizer_int_chain_out1(\alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.altera_reset_synchronizer_int_chain_1(altera_reset_synchronizer_int_chain_1),
	.clk(clk_clk));

nios_mcu_altera_reset_synchronizer_1 alt_rst_sync_uq1(
	.altera_reset_synchronizer_int_chain_out1(\alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.clk(clk_clk),
	.reset_reset_n(reset_reset_n));

dffeas r_sync_rst(
	.clk(clk_clk),
	.d(\WideOr0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_sync_rst1),
	.prn(vcc));
defparam r_sync_rst.is_wysiwyg = "true";
defparam r_sync_rst.power_up = "low";

dffeas r_early_rst(
	.clk(clk_clk),
	.d(\always2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_early_rst1),
	.prn(vcc));
defparam r_early_rst.is_wysiwyg = "true";
defparam r_early_rst.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk_clk),
	.d(\alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[2] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[2]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[2] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[2] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[3] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[3]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[3] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[3] .power_up = "low";

cycloneive_lcell_comb \altera_reset_synchronizer_int_chain[4]~0 (
	.dataa(\altera_reset_synchronizer_int_chain[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\altera_reset_synchronizer_int_chain[4]~0_combout ),
	.cout());
defparam \altera_reset_synchronizer_int_chain[4]~0 .lut_mask = 16'h5555;
defparam \altera_reset_synchronizer_int_chain[4]~0 .sum_lutc_input = "datac";

dffeas \altera_reset_synchronizer_int_chain[4] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[4]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[4]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[4] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[4] .power_up = "low";

dffeas \r_sync_rst_chain[3] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[3]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[3] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[3] .power_up = "low";

cycloneive_lcell_comb \r_sync_rst_chain~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\altera_reset_synchronizer_int_chain[2]~q ),
	.datad(\r_sync_rst_chain[3]~q ),
	.cin(gnd),
	.combout(\r_sync_rst_chain~1_combout ),
	.cout());
defparam \r_sync_rst_chain~1 .lut_mask = 16'hFFF0;
defparam \r_sync_rst_chain~1 .sum_lutc_input = "datac";

dffeas \r_sync_rst_chain[2] (
	.clk(clk_clk),
	.d(\r_sync_rst_chain~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[2]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[2] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[2] .power_up = "low";

cycloneive_lcell_comb \r_sync_rst_chain~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\altera_reset_synchronizer_int_chain[2]~q ),
	.datad(\r_sync_rst_chain[2]~q ),
	.cin(gnd),
	.combout(\r_sync_rst_chain~0_combout ),
	.cout());
defparam \r_sync_rst_chain~0 .lut_mask = 16'hFFF0;
defparam \r_sync_rst_chain~0 .sum_lutc_input = "datac";

dffeas \r_sync_rst_chain[1] (
	.clk(clk_clk),
	.d(\r_sync_rst_chain~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[1]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[1] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[1] .power_up = "low";

cycloneive_lcell_comb \WideOr0~0 (
	.dataa(\altera_reset_synchronizer_int_chain[4]~q ),
	.datab(r_sync_rst1),
	.datac(gnd),
	.datad(\r_sync_rst_chain[1]~q ),
	.cin(gnd),
	.combout(\WideOr0~0_combout ),
	.cout());
defparam \WideOr0~0 .lut_mask = 16'hEEFF;
defparam \WideOr0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always2~0 (
	.dataa(\alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\r_sync_rst_chain[2]~q ),
	.cin(gnd),
	.combout(\always2~0_combout ),
	.cout());
defparam \always2~0 .lut_mask = 16'hAAFF;
defparam \always2~0 .sum_lutc_input = "datac";

endmodule

module nios_mcu_altera_reset_synchronizer (
	altera_reset_synchronizer_int_chain_out1,
	altera_reset_synchronizer_int_chain_1,
	clk)/* synthesis synthesis_greybox=1 */;
output 	altera_reset_synchronizer_int_chain_out1;
output 	altera_reset_synchronizer_int_chain_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

cycloneive_lcell_comb \altera_reset_synchronizer_int_chain[1]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(altera_reset_synchronizer_int_chain_1),
	.cout());
defparam \altera_reset_synchronizer_int_chain[1]~0 .lut_mask = 16'h0000;
defparam \altera_reset_synchronizer_int_chain[1]~0 .sum_lutc_input = "datac";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(altera_reset_synchronizer_int_chain_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module nios_mcu_altera_reset_synchronizer_1 (
	altera_reset_synchronizer_int_chain_out1,
	clk,
	reset_reset_n)/* synthesis synthesis_greybox=1 */;
output 	altera_reset_synchronizer_int_chain_out1;
input 	clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module nios_mcu_AvalonSlave (
	W_alu_result_3,
	W_alu_result_2,
	d_writedata_24,
	d_writedata_25,
	d_writedata_26,
	d_writedata_27,
	d_writedata_28,
	d_writedata_29,
	d_writedata_30,
	d_writedata_31,
	d_writedata_0,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	m0_write,
	Equal2,
	dRead1,
	m0_read,
	Read,
	sReadCountPipelined_0,
	Equal21,
	ReadData_0,
	d_byteenable_0,
	d_writedata_22,
	d_byteenable_2,
	d_writedata_23,
	d_byteenable_3,
	d_writedata_11,
	d_byteenable_1,
	d_writedata_13,
	d_writedata_16,
	d_writedata_12,
	d_writedata_14,
	d_writedata_15,
	d_writedata_18,
	d_writedata_17,
	d_writedata_10,
	d_writedata_9,
	d_writedata_8,
	d_writedata_21,
	d_writedata_19,
	d_writedata_20,
	ReadData_1,
	ReadData_2,
	ReadData_3,
	ReadData_4,
	ReadData_5,
	ReadData_6,
	ReadData_7,
	ReadData_8,
	ReadData_12,
	ReadData_11,
	ReadData_10,
	ReadData_9,
	ReadData_15,
	ReadData_14,
	ReadData_13,
	ReadData_16,
	ReadData_20,
	ReadData_19,
	ReadData_18,
	ReadData_17,
	ReadData_23,
	ReadData_22,
	ReadData_21,
	ReadData_24,
	ReadData_31,
	ReadData_30,
	ReadData_29,
	ReadData_28,
	ReadData_27,
	ReadData_26,
	ReadData_25,
	Clk,
	Reset)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_3;
input 	W_alu_result_2;
input 	d_writedata_24;
input 	d_writedata_25;
input 	d_writedata_26;
input 	d_writedata_27;
input 	d_writedata_28;
input 	d_writedata_29;
input 	d_writedata_30;
input 	d_writedata_31;
input 	d_writedata_0;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	d_writedata_6;
input 	d_writedata_7;
input 	m0_write;
input 	Equal2;
output 	dRead1;
input 	m0_read;
input 	Read;
output 	sReadCountPipelined_0;
output 	Equal21;
output 	ReadData_0;
input 	d_byteenable_0;
input 	d_writedata_22;
input 	d_byteenable_2;
input 	d_writedata_23;
input 	d_byteenable_3;
input 	d_writedata_11;
input 	d_byteenable_1;
input 	d_writedata_13;
input 	d_writedata_16;
input 	d_writedata_12;
input 	d_writedata_14;
input 	d_writedata_15;
input 	d_writedata_18;
input 	d_writedata_17;
input 	d_writedata_10;
input 	d_writedata_9;
input 	d_writedata_8;
input 	d_writedata_21;
input 	d_writedata_19;
input 	d_writedata_20;
output 	ReadData_1;
output 	ReadData_2;
output 	ReadData_3;
output 	ReadData_4;
output 	ReadData_5;
output 	ReadData_6;
output 	ReadData_7;
output 	ReadData_8;
output 	ReadData_12;
output 	ReadData_11;
output 	ReadData_10;
output 	ReadData_9;
output 	ReadData_15;
output 	ReadData_14;
output 	ReadData_13;
output 	ReadData_16;
output 	ReadData_20;
output 	ReadData_19;
output 	ReadData_18;
output 	ReadData_17;
output 	ReadData_23;
output 	ReadData_22;
output 	ReadData_21;
output 	ReadData_24;
output 	ReadData_31;
output 	ReadData_30;
output 	ReadData_29;
output 	ReadData_28;
output 	ReadData_27;
output 	ReadData_26;
output 	ReadData_25;
input 	Clk;
input 	Reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \sRegByteEnable[24]~0_combout ;
wire \sRegByteEnable[24]~1_combout ;
wire \sRegByteEnable[0]~2_combout ;
wire \sRegByteEnable[0]~q ;
wire \sReadCount[0]~32_combout ;
wire \sReadCount[0]~34_combout ;
wire \sReadCount[0]~q ;
wire \Mux31~0_combout ;
wire \sReg[0]~0_combout ;
wire \sReg[0]~q ;
wire \ReadData[0]~0_combout ;
wire \sReadCountPipelined[0]~33_combout ;
wire \sReadCountPipelined[0]~q ;
wire \sReadCount[0]~33 ;
wire \sReadCount[1]~35_combout ;
wire \sReadCount[1]~q ;
wire \sRegByteEnable[1]~q ;
wire \sReg[1]~q ;
wire \ReadData[1]~2_combout ;
wire \sReadCountPipelined[0]~34 ;
wire \sReadCountPipelined[1]~35_combout ;
wire \sReadCountPipelined[1]~q ;
wire \sRegByteEnable[2]~q ;
wire \sReadCount[1]~36 ;
wire \sReadCount[2]~37_combout ;
wire \sReadCount[2]~q ;
wire \sReg[2]~q ;
wire \ReadData[2]~4_combout ;
wire \sReadCountPipelined[1]~36 ;
wire \sReadCountPipelined[2]~37_combout ;
wire \sReadCountPipelined[2]~q ;
wire \sReadCount[2]~38 ;
wire \sReadCount[3]~39_combout ;
wire \sReadCount[3]~q ;
wire \sRegByteEnable[3]~q ;
wire \sReg[3]~q ;
wire \ReadData[3]~6_combout ;
wire \sReadCountPipelined[2]~38 ;
wire \sReadCountPipelined[3]~39_combout ;
wire \sReadCountPipelined[3]~q ;
wire \sRegByteEnable[4]~q ;
wire \sReadCount[3]~40 ;
wire \sReadCount[4]~41_combout ;
wire \sReadCount[4]~q ;
wire \sReg[4]~q ;
wire \ReadData[4]~8_combout ;
wire \sReadCountPipelined[3]~40 ;
wire \sReadCountPipelined[4]~41_combout ;
wire \sReadCountPipelined[4]~q ;
wire \sReadCount[4]~42 ;
wire \sReadCount[5]~43_combout ;
wire \sReadCount[5]~q ;
wire \sRegByteEnable[5]~q ;
wire \sReg[5]~q ;
wire \ReadData[5]~10_combout ;
wire \sReadCountPipelined[4]~42 ;
wire \sReadCountPipelined[5]~43_combout ;
wire \sReadCountPipelined[5]~q ;
wire \sRegByteEnable[6]~q ;
wire \sReadCount[5]~44 ;
wire \sReadCount[6]~45_combout ;
wire \sReadCount[6]~q ;
wire \sReg[6]~q ;
wire \ReadData[6]~12_combout ;
wire \sReadCountPipelined[5]~44 ;
wire \sReadCountPipelined[6]~45_combout ;
wire \sReadCountPipelined[6]~q ;
wire \sReadCount[6]~46 ;
wire \sReadCount[7]~47_combout ;
wire \sReadCount[7]~q ;
wire \sRegByteEnable[7]~q ;
wire \sReg[7]~q ;
wire \ReadData[7]~14_combout ;
wire \sReadCountPipelined[6]~46 ;
wire \sReadCountPipelined[7]~47_combout ;
wire \sReadCountPipelined[7]~q ;
wire \sRegByteEnable[8]~3_combout ;
wire \sRegByteEnable[8]~q ;
wire \sReadCount[7]~48 ;
wire \sReadCount[8]~49_combout ;
wire \sReadCount[8]~q ;
wire \sReg[8]~q ;
wire \ReadData[8]~16_combout ;
wire \sReadCountPipelined[7]~48 ;
wire \sReadCountPipelined[8]~49_combout ;
wire \sReadCountPipelined[8]~q ;
wire \sRegByteEnable[12]~q ;
wire \sReadCount[8]~50 ;
wire \sReadCount[9]~51_combout ;
wire \sReadCount[9]~q ;
wire \sReadCount[9]~52 ;
wire \sReadCount[10]~53_combout ;
wire \sReadCount[10]~q ;
wire \sReadCount[10]~54 ;
wire \sReadCount[11]~55_combout ;
wire \sReadCount[11]~q ;
wire \sReadCount[11]~56 ;
wire \sReadCount[12]~57_combout ;
wire \sReadCount[12]~q ;
wire \sReg[12]~q ;
wire \ReadData[12]~18_combout ;
wire \sReadCountPipelined[8]~50 ;
wire \sReadCountPipelined[9]~51_combout ;
wire \sReadCountPipelined[9]~q ;
wire \sReadCountPipelined[9]~52 ;
wire \sReadCountPipelined[10]~53_combout ;
wire \sReadCountPipelined[10]~q ;
wire \sReadCountPipelined[10]~54 ;
wire \sReadCountPipelined[11]~55_combout ;
wire \sReadCountPipelined[11]~q ;
wire \sReadCountPipelined[11]~56 ;
wire \sReadCountPipelined[12]~57_combout ;
wire \sReadCountPipelined[12]~q ;
wire \sRegByteEnable[11]~q ;
wire \sReg[11]~q ;
wire \ReadData[11]~20_combout ;
wire \sRegByteEnable[10]~q ;
wire \sReg[10]~q ;
wire \ReadData[10]~22_combout ;
wire \sRegByteEnable[9]~q ;
wire \sReg[9]~q ;
wire \ReadData[9]~24_combout ;
wire \sReadCount[12]~58 ;
wire \sReadCount[13]~59_combout ;
wire \sReadCount[13]~q ;
wire \sReadCount[13]~60 ;
wire \sReadCount[14]~61_combout ;
wire \sReadCount[14]~q ;
wire \sReadCount[14]~62 ;
wire \sReadCount[15]~63_combout ;
wire \sReadCount[15]~q ;
wire \sRegByteEnable[15]~q ;
wire \sReg[15]~q ;
wire \ReadData[15]~26_combout ;
wire \sReadCountPipelined[12]~58 ;
wire \sReadCountPipelined[13]~59_combout ;
wire \sReadCountPipelined[13]~q ;
wire \sReadCountPipelined[13]~60 ;
wire \sReadCountPipelined[14]~61_combout ;
wire \sReadCountPipelined[14]~q ;
wire \sReadCountPipelined[14]~62 ;
wire \sReadCountPipelined[15]~63_combout ;
wire \sReadCountPipelined[15]~q ;
wire \sRegByteEnable[14]~q ;
wire \sReg[14]~q ;
wire \ReadData[14]~28_combout ;
wire \sRegByteEnable[13]~q ;
wire \sReg[13]~q ;
wire \ReadData[13]~30_combout ;
wire \sRegByteEnable[16]~4_combout ;
wire \sRegByteEnable[16]~q ;
wire \sReadCount[15]~64 ;
wire \sReadCount[16]~65_combout ;
wire \sReadCount[16]~q ;
wire \sReg[16]~q ;
wire \ReadData[16]~32_combout ;
wire \sReadCountPipelined[15]~64 ;
wire \sReadCountPipelined[16]~65_combout ;
wire \sReadCountPipelined[16]~q ;
wire \sRegByteEnable[20]~q ;
wire \sReadCount[16]~66 ;
wire \sReadCount[17]~67_combout ;
wire \sReadCount[17]~q ;
wire \sReadCount[17]~68 ;
wire \sReadCount[18]~69_combout ;
wire \sReadCount[18]~q ;
wire \sReadCount[18]~70 ;
wire \sReadCount[19]~71_combout ;
wire \sReadCount[19]~q ;
wire \sReadCount[19]~72 ;
wire \sReadCount[20]~73_combout ;
wire \sReadCount[20]~q ;
wire \sReg[20]~q ;
wire \ReadData[20]~34_combout ;
wire \sReadCountPipelined[16]~66 ;
wire \sReadCountPipelined[17]~67_combout ;
wire \sReadCountPipelined[17]~q ;
wire \sReadCountPipelined[17]~68 ;
wire \sReadCountPipelined[18]~69_combout ;
wire \sReadCountPipelined[18]~q ;
wire \sReadCountPipelined[18]~70 ;
wire \sReadCountPipelined[19]~71_combout ;
wire \sReadCountPipelined[19]~q ;
wire \sReadCountPipelined[19]~72 ;
wire \sReadCountPipelined[20]~73_combout ;
wire \sReadCountPipelined[20]~q ;
wire \sRegByteEnable[19]~q ;
wire \sReg[19]~q ;
wire \ReadData[19]~36_combout ;
wire \sRegByteEnable[18]~q ;
wire \sReg[18]~q ;
wire \ReadData[18]~38_combout ;
wire \sRegByteEnable[17]~q ;
wire \sReg[17]~q ;
wire \ReadData[17]~40_combout ;
wire \sReadCount[20]~74 ;
wire \sReadCount[21]~75_combout ;
wire \sReadCount[21]~q ;
wire \sReadCount[21]~76 ;
wire \sReadCount[22]~77_combout ;
wire \sReadCount[22]~q ;
wire \sReadCount[22]~78 ;
wire \sReadCount[23]~79_combout ;
wire \sReadCount[23]~q ;
wire \sRegByteEnable[23]~q ;
wire \sReg[23]~q ;
wire \ReadData[23]~42_combout ;
wire \sReadCountPipelined[20]~74 ;
wire \sReadCountPipelined[21]~75_combout ;
wire \sReadCountPipelined[21]~q ;
wire \sReadCountPipelined[21]~76 ;
wire \sReadCountPipelined[22]~77_combout ;
wire \sReadCountPipelined[22]~q ;
wire \sReadCountPipelined[22]~78 ;
wire \sReadCountPipelined[23]~79_combout ;
wire \sReadCountPipelined[23]~q ;
wire \sRegByteEnable[22]~q ;
wire \sReg[22]~q ;
wire \ReadData[22]~44_combout ;
wire \sRegByteEnable[21]~q ;
wire \sReg[21]~q ;
wire \ReadData[21]~46_combout ;
wire \sRegByteEnable[24]~5_combout ;
wire \sRegByteEnable[24]~q ;
wire \sReadCount[23]~80 ;
wire \sReadCount[24]~81_combout ;
wire \sReadCount[24]~q ;
wire \sReg[24]~q ;
wire \ReadData[24]~48_combout ;
wire \sReadCountPipelined[23]~80 ;
wire \sReadCountPipelined[24]~81_combout ;
wire \sReadCountPipelined[24]~q ;
wire \sReadCount[24]~82 ;
wire \sReadCount[25]~83_combout ;
wire \sReadCount[25]~q ;
wire \sReadCount[25]~84 ;
wire \sReadCount[26]~85_combout ;
wire \sReadCount[26]~q ;
wire \sReadCount[26]~86 ;
wire \sReadCount[27]~87_combout ;
wire \sReadCount[27]~q ;
wire \sReadCount[27]~88 ;
wire \sReadCount[28]~89_combout ;
wire \sReadCount[28]~q ;
wire \sReadCount[28]~90 ;
wire \sReadCount[29]~91_combout ;
wire \sReadCount[29]~q ;
wire \sReadCount[29]~92 ;
wire \sReadCount[30]~93_combout ;
wire \sReadCount[30]~q ;
wire \sReadCount[30]~94 ;
wire \sReadCount[31]~95_combout ;
wire \sReadCount[31]~q ;
wire \sRegByteEnable[31]~q ;
wire \sReg[31]~q ;
wire \ReadData[31]~50_combout ;
wire \sReadCountPipelined[24]~82 ;
wire \sReadCountPipelined[25]~83_combout ;
wire \sReadCountPipelined[25]~q ;
wire \sReadCountPipelined[25]~84 ;
wire \sReadCountPipelined[26]~85_combout ;
wire \sReadCountPipelined[26]~q ;
wire \sReadCountPipelined[26]~86 ;
wire \sReadCountPipelined[27]~87_combout ;
wire \sReadCountPipelined[27]~q ;
wire \sReadCountPipelined[27]~88 ;
wire \sReadCountPipelined[28]~89_combout ;
wire \sReadCountPipelined[28]~q ;
wire \sReadCountPipelined[28]~90 ;
wire \sReadCountPipelined[29]~91_combout ;
wire \sReadCountPipelined[29]~q ;
wire \sReadCountPipelined[29]~92 ;
wire \sReadCountPipelined[30]~93_combout ;
wire \sReadCountPipelined[30]~q ;
wire \sReadCountPipelined[30]~94 ;
wire \sReadCountPipelined[31]~95_combout ;
wire \sReadCountPipelined[31]~q ;
wire \sRegByteEnable[30]~q ;
wire \sReg[30]~q ;
wire \ReadData[30]~52_combout ;
wire \sRegByteEnable[29]~q ;
wire \sReg[29]~q ;
wire \ReadData[29]~54_combout ;
wire \sRegByteEnable[28]~q ;
wire \sReg[28]~q ;
wire \ReadData[28]~56_combout ;
wire \sRegByteEnable[27]~q ;
wire \sReg[27]~q ;
wire \ReadData[27]~58_combout ;
wire \sRegByteEnable[26]~q ;
wire \sReg[26]~q ;
wire \ReadData[26]~60_combout ;
wire \sRegByteEnable[25]~q ;
wire \sReg[25]~q ;
wire \ReadData[25]~62_combout ;


dffeas dRead(
	.clk(Clk),
	.d(Read),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dRead1),
	.prn(vcc));
defparam dRead.is_wysiwyg = "true";
defparam dRead.power_up = "low";

cycloneive_lcell_comb \sReadCountPipelined[0]~32 (
	.dataa(W_alu_result_3),
	.datab(W_alu_result_2),
	.datac(Read),
	.datad(gnd),
	.cin(gnd),
	.combout(sReadCountPipelined_0),
	.cout());
defparam \sReadCountPipelined[0]~32 .lut_mask = 16'hFEFE;
defparam \sReadCountPipelined[0]~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal2~0 (
	.dataa(W_alu_result_3),
	.datab(W_alu_result_2),
	.datac(Read),
	.datad(dRead1),
	.cin(gnd),
	.combout(Equal21),
	.cout());
defparam \Equal2~0 .lut_mask = 16'hFEFF;
defparam \Equal2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ReadData[0]~1 (
	.dataa(\sRegByteEnable[0]~q ),
	.datab(W_alu_result_2),
	.datac(\ReadData[0]~0_combout ),
	.datad(\sReadCountPipelined[0]~q ),
	.cin(gnd),
	.combout(ReadData_0),
	.cout());
defparam \ReadData[0]~1 .lut_mask = 16'hFFBE;
defparam \ReadData[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ReadData[1]~3 (
	.dataa(\sReadCount[1]~q ),
	.datab(W_alu_result_3),
	.datac(\ReadData[1]~2_combout ),
	.datad(\sReadCountPipelined[1]~q ),
	.cin(gnd),
	.combout(ReadData_1),
	.cout());
defparam \ReadData[1]~3 .lut_mask = 16'hFFBE;
defparam \ReadData[1]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ReadData[2]~5 (
	.dataa(\sRegByteEnable[2]~q ),
	.datab(W_alu_result_2),
	.datac(\ReadData[2]~4_combout ),
	.datad(\sReadCountPipelined[2]~q ),
	.cin(gnd),
	.combout(ReadData_2),
	.cout());
defparam \ReadData[2]~5 .lut_mask = 16'hFFBE;
defparam \ReadData[2]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ReadData[3]~7 (
	.dataa(\sReadCount[3]~q ),
	.datab(W_alu_result_3),
	.datac(\ReadData[3]~6_combout ),
	.datad(\sReadCountPipelined[3]~q ),
	.cin(gnd),
	.combout(ReadData_3),
	.cout());
defparam \ReadData[3]~7 .lut_mask = 16'hFFBE;
defparam \ReadData[3]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ReadData[4]~9 (
	.dataa(\sRegByteEnable[4]~q ),
	.datab(W_alu_result_2),
	.datac(\ReadData[4]~8_combout ),
	.datad(\sReadCountPipelined[4]~q ),
	.cin(gnd),
	.combout(ReadData_4),
	.cout());
defparam \ReadData[4]~9 .lut_mask = 16'hFFBE;
defparam \ReadData[4]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ReadData[5]~11 (
	.dataa(\sReadCount[5]~q ),
	.datab(W_alu_result_3),
	.datac(\ReadData[5]~10_combout ),
	.datad(\sReadCountPipelined[5]~q ),
	.cin(gnd),
	.combout(ReadData_5),
	.cout());
defparam \ReadData[5]~11 .lut_mask = 16'hFFBE;
defparam \ReadData[5]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ReadData[6]~13 (
	.dataa(\sRegByteEnable[6]~q ),
	.datab(W_alu_result_2),
	.datac(\ReadData[6]~12_combout ),
	.datad(\sReadCountPipelined[6]~q ),
	.cin(gnd),
	.combout(ReadData_6),
	.cout());
defparam \ReadData[6]~13 .lut_mask = 16'hFFBE;
defparam \ReadData[6]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ReadData[7]~15 (
	.dataa(\sReadCount[7]~q ),
	.datab(W_alu_result_3),
	.datac(\ReadData[7]~14_combout ),
	.datad(\sReadCountPipelined[7]~q ),
	.cin(gnd),
	.combout(ReadData_7),
	.cout());
defparam \ReadData[7]~15 .lut_mask = 16'hFFBE;
defparam \ReadData[7]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ReadData[8]~17 (
	.dataa(\sRegByteEnable[8]~q ),
	.datab(W_alu_result_2),
	.datac(\ReadData[8]~16_combout ),
	.datad(\sReadCountPipelined[8]~q ),
	.cin(gnd),
	.combout(ReadData_8),
	.cout());
defparam \ReadData[8]~17 .lut_mask = 16'hFFBE;
defparam \ReadData[8]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ReadData[12]~19 (
	.dataa(\sRegByteEnable[12]~q ),
	.datab(W_alu_result_2),
	.datac(\ReadData[12]~18_combout ),
	.datad(\sReadCountPipelined[12]~q ),
	.cin(gnd),
	.combout(ReadData_12),
	.cout());
defparam \ReadData[12]~19 .lut_mask = 16'hFFBE;
defparam \ReadData[12]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ReadData[11]~21 (
	.dataa(\sReadCount[11]~q ),
	.datab(W_alu_result_3),
	.datac(\ReadData[11]~20_combout ),
	.datad(\sReadCountPipelined[11]~q ),
	.cin(gnd),
	.combout(ReadData_11),
	.cout());
defparam \ReadData[11]~21 .lut_mask = 16'hFFBE;
defparam \ReadData[11]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ReadData[10]~23 (
	.dataa(\sRegByteEnable[10]~q ),
	.datab(W_alu_result_2),
	.datac(\ReadData[10]~22_combout ),
	.datad(\sReadCountPipelined[10]~q ),
	.cin(gnd),
	.combout(ReadData_10),
	.cout());
defparam \ReadData[10]~23 .lut_mask = 16'hFFBE;
defparam \ReadData[10]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ReadData[9]~25 (
	.dataa(\sReadCount[9]~q ),
	.datab(W_alu_result_3),
	.datac(\ReadData[9]~24_combout ),
	.datad(\sReadCountPipelined[9]~q ),
	.cin(gnd),
	.combout(ReadData_9),
	.cout());
defparam \ReadData[9]~25 .lut_mask = 16'hFFBE;
defparam \ReadData[9]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ReadData[15]~27 (
	.dataa(\sReadCount[15]~q ),
	.datab(W_alu_result_3),
	.datac(\ReadData[15]~26_combout ),
	.datad(\sReadCountPipelined[15]~q ),
	.cin(gnd),
	.combout(ReadData_15),
	.cout());
defparam \ReadData[15]~27 .lut_mask = 16'hFFBE;
defparam \ReadData[15]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ReadData[14]~29 (
	.dataa(\sRegByteEnable[14]~q ),
	.datab(W_alu_result_2),
	.datac(\ReadData[14]~28_combout ),
	.datad(\sReadCountPipelined[14]~q ),
	.cin(gnd),
	.combout(ReadData_14),
	.cout());
defparam \ReadData[14]~29 .lut_mask = 16'hFFBE;
defparam \ReadData[14]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ReadData[13]~31 (
	.dataa(\sReadCount[13]~q ),
	.datab(W_alu_result_3),
	.datac(\ReadData[13]~30_combout ),
	.datad(\sReadCountPipelined[13]~q ),
	.cin(gnd),
	.combout(ReadData_13),
	.cout());
defparam \ReadData[13]~31 .lut_mask = 16'hFFBE;
defparam \ReadData[13]~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ReadData[16]~33 (
	.dataa(\sRegByteEnable[16]~q ),
	.datab(W_alu_result_2),
	.datac(\ReadData[16]~32_combout ),
	.datad(\sReadCountPipelined[16]~q ),
	.cin(gnd),
	.combout(ReadData_16),
	.cout());
defparam \ReadData[16]~33 .lut_mask = 16'hFFBE;
defparam \ReadData[16]~33 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ReadData[20]~35 (
	.dataa(\sRegByteEnable[20]~q ),
	.datab(W_alu_result_2),
	.datac(\ReadData[20]~34_combout ),
	.datad(\sReadCountPipelined[20]~q ),
	.cin(gnd),
	.combout(ReadData_20),
	.cout());
defparam \ReadData[20]~35 .lut_mask = 16'hFFBE;
defparam \ReadData[20]~35 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ReadData[19]~37 (
	.dataa(\sReadCount[19]~q ),
	.datab(W_alu_result_3),
	.datac(\ReadData[19]~36_combout ),
	.datad(\sReadCountPipelined[19]~q ),
	.cin(gnd),
	.combout(ReadData_19),
	.cout());
defparam \ReadData[19]~37 .lut_mask = 16'hFFBE;
defparam \ReadData[19]~37 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ReadData[18]~39 (
	.dataa(\sRegByteEnable[18]~q ),
	.datab(W_alu_result_2),
	.datac(\ReadData[18]~38_combout ),
	.datad(\sReadCountPipelined[18]~q ),
	.cin(gnd),
	.combout(ReadData_18),
	.cout());
defparam \ReadData[18]~39 .lut_mask = 16'hFFBE;
defparam \ReadData[18]~39 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ReadData[17]~41 (
	.dataa(\sReadCount[17]~q ),
	.datab(W_alu_result_3),
	.datac(\ReadData[17]~40_combout ),
	.datad(\sReadCountPipelined[17]~q ),
	.cin(gnd),
	.combout(ReadData_17),
	.cout());
defparam \ReadData[17]~41 .lut_mask = 16'hFFBE;
defparam \ReadData[17]~41 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ReadData[23]~43 (
	.dataa(\sReadCount[23]~q ),
	.datab(W_alu_result_3),
	.datac(\ReadData[23]~42_combout ),
	.datad(\sReadCountPipelined[23]~q ),
	.cin(gnd),
	.combout(ReadData_23),
	.cout());
defparam \ReadData[23]~43 .lut_mask = 16'hFFBE;
defparam \ReadData[23]~43 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ReadData[22]~45 (
	.dataa(\sRegByteEnable[22]~q ),
	.datab(W_alu_result_2),
	.datac(\ReadData[22]~44_combout ),
	.datad(\sReadCountPipelined[22]~q ),
	.cin(gnd),
	.combout(ReadData_22),
	.cout());
defparam \ReadData[22]~45 .lut_mask = 16'hFFBE;
defparam \ReadData[22]~45 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ReadData[21]~47 (
	.dataa(\sReadCount[21]~q ),
	.datab(W_alu_result_3),
	.datac(\ReadData[21]~46_combout ),
	.datad(\sReadCountPipelined[21]~q ),
	.cin(gnd),
	.combout(ReadData_21),
	.cout());
defparam \ReadData[21]~47 .lut_mask = 16'hFFBE;
defparam \ReadData[21]~47 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ReadData[24]~49 (
	.dataa(\sRegByteEnable[24]~q ),
	.datab(W_alu_result_2),
	.datac(\ReadData[24]~48_combout ),
	.datad(\sReadCountPipelined[24]~q ),
	.cin(gnd),
	.combout(ReadData_24),
	.cout());
defparam \ReadData[24]~49 .lut_mask = 16'hFFBE;
defparam \ReadData[24]~49 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ReadData[31]~51 (
	.dataa(\sReadCount[31]~q ),
	.datab(W_alu_result_3),
	.datac(\ReadData[31]~50_combout ),
	.datad(\sReadCountPipelined[31]~q ),
	.cin(gnd),
	.combout(ReadData_31),
	.cout());
defparam \ReadData[31]~51 .lut_mask = 16'hFFBE;
defparam \ReadData[31]~51 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ReadData[30]~53 (
	.dataa(\sRegByteEnable[30]~q ),
	.datab(W_alu_result_2),
	.datac(\ReadData[30]~52_combout ),
	.datad(\sReadCountPipelined[30]~q ),
	.cin(gnd),
	.combout(ReadData_30),
	.cout());
defparam \ReadData[30]~53 .lut_mask = 16'hFFBE;
defparam \ReadData[30]~53 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ReadData[29]~55 (
	.dataa(\sReadCount[29]~q ),
	.datab(W_alu_result_3),
	.datac(\ReadData[29]~54_combout ),
	.datad(\sReadCountPipelined[29]~q ),
	.cin(gnd),
	.combout(ReadData_29),
	.cout());
defparam \ReadData[29]~55 .lut_mask = 16'hFFBE;
defparam \ReadData[29]~55 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ReadData[28]~57 (
	.dataa(\sRegByteEnable[28]~q ),
	.datab(W_alu_result_2),
	.datac(\ReadData[28]~56_combout ),
	.datad(\sReadCountPipelined[28]~q ),
	.cin(gnd),
	.combout(ReadData_28),
	.cout());
defparam \ReadData[28]~57 .lut_mask = 16'hFFBE;
defparam \ReadData[28]~57 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ReadData[27]~59 (
	.dataa(\sReadCount[27]~q ),
	.datab(W_alu_result_3),
	.datac(\ReadData[27]~58_combout ),
	.datad(\sReadCountPipelined[27]~q ),
	.cin(gnd),
	.combout(ReadData_27),
	.cout());
defparam \ReadData[27]~59 .lut_mask = 16'hFFBE;
defparam \ReadData[27]~59 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ReadData[26]~61 (
	.dataa(\sRegByteEnable[26]~q ),
	.datab(W_alu_result_2),
	.datac(\ReadData[26]~60_combout ),
	.datad(\sReadCountPipelined[26]~q ),
	.cin(gnd),
	.combout(ReadData_26),
	.cout());
defparam \ReadData[26]~61 .lut_mask = 16'hFFBE;
defparam \ReadData[26]~61 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ReadData[25]~63 (
	.dataa(\sReadCount[25]~q ),
	.datab(W_alu_result_3),
	.datac(\ReadData[25]~62_combout ),
	.datad(\sReadCountPipelined[25]~q ),
	.cin(gnd),
	.combout(ReadData_25),
	.cout());
defparam \ReadData[25]~63 .lut_mask = 16'hFFBE;
defparam \ReadData[25]~63 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sRegByteEnable[24]~0 (
	.dataa(W_alu_result_2),
	.datab(Reset),
	.datac(gnd),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(\sRegByteEnable[24]~0_combout ),
	.cout());
defparam \sRegByteEnable[24]~0 .lut_mask = 16'hEEFF;
defparam \sRegByteEnable[24]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sRegByteEnable[24]~1 (
	.dataa(m0_write),
	.datab(Equal2),
	.datac(m0_read),
	.datad(\sRegByteEnable[24]~0_combout ),
	.cin(gnd),
	.combout(\sRegByteEnable[24]~1_combout ),
	.cout());
defparam \sRegByteEnable[24]~1 .lut_mask = 16'hFFFE;
defparam \sRegByteEnable[24]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sRegByteEnable[0]~2 (
	.dataa(d_byteenable_0),
	.datab(\sRegByteEnable[24]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sRegByteEnable[0]~2_combout ),
	.cout());
defparam \sRegByteEnable[0]~2 .lut_mask = 16'hEEEE;
defparam \sRegByteEnable[0]~2 .sum_lutc_input = "datac";

dffeas \sRegByteEnable[0] (
	.clk(Clk),
	.d(d_writedata_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sRegByteEnable[0]~2_combout ),
	.q(\sRegByteEnable[0]~q ),
	.prn(vcc));
defparam \sRegByteEnable[0] .is_wysiwyg = "true";
defparam \sRegByteEnable[0] .power_up = "low";

cycloneive_lcell_comb \sReadCount[0]~32 (
	.dataa(\sReadCount[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\sReadCount[0]~32_combout ),
	.cout(\sReadCount[0]~33 ));
defparam \sReadCount[0]~32 .lut_mask = 16'h55AA;
defparam \sReadCount[0]~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sReadCount[0]~34 (
	.dataa(W_alu_result_3),
	.datab(Read),
	.datac(gnd),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\sReadCount[0]~34_combout ),
	.cout());
defparam \sReadCount[0]~34 .lut_mask = 16'hEEFF;
defparam \sReadCount[0]~34 .sum_lutc_input = "datac";

dffeas \sReadCount[0] (
	.clk(Clk),
	.d(\sReadCount[0]~32_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReadCount[0]~34_combout ),
	.q(\sReadCount[0]~q ),
	.prn(vcc));
defparam \sReadCount[0] .is_wysiwyg = "true";
defparam \sReadCount[0] .power_up = "low";

cycloneive_lcell_comb \Mux31~0 (
	.dataa(W_alu_result_3),
	.datab(W_alu_result_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux31~0_combout ),
	.cout());
defparam \Mux31~0 .lut_mask = 16'hEEEE;
defparam \Mux31~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sReg[0]~0 (
	.dataa(m0_write),
	.datab(Equal2),
	.datac(m0_read),
	.datad(\Mux31~0_combout ),
	.cin(gnd),
	.combout(\sReg[0]~0_combout ),
	.cout());
defparam \sReg[0]~0 .lut_mask = 16'hFEFF;
defparam \sReg[0]~0 .sum_lutc_input = "datac";

dffeas \sReg[0] (
	.clk(Clk),
	.d(d_writedata_0),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReg[0]~0_combout ),
	.q(\sReg[0]~q ),
	.prn(vcc));
defparam \sReg[0] .is_wysiwyg = "true";
defparam \sReg[0] .power_up = "low";

cycloneive_lcell_comb \ReadData[0]~0 (
	.dataa(W_alu_result_2),
	.datab(\sReadCount[0]~q ),
	.datac(W_alu_result_3),
	.datad(\sReg[0]~q ),
	.cin(gnd),
	.combout(\ReadData[0]~0_combout ),
	.cout());
defparam \ReadData[0]~0 .lut_mask = 16'hFFDE;
defparam \ReadData[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sReadCountPipelined[0]~33 (
	.dataa(dRead1),
	.datab(\sReadCountPipelined[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\sReadCountPipelined[0]~33_combout ),
	.cout(\sReadCountPipelined[0]~34 ));
defparam \sReadCountPipelined[0]~33 .lut_mask = 16'h66DD;
defparam \sReadCountPipelined[0]~33 .sum_lutc_input = "datac";

dffeas \sReadCountPipelined[0] (
	.clk(Clk),
	.d(\sReadCountPipelined[0]~33_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sReadCountPipelined_0),
	.q(\sReadCountPipelined[0]~q ),
	.prn(vcc));
defparam \sReadCountPipelined[0] .is_wysiwyg = "true";
defparam \sReadCountPipelined[0] .power_up = "low";

cycloneive_lcell_comb \sReadCount[1]~35 (
	.dataa(\sReadCount[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCount[0]~33 ),
	.combout(\sReadCount[1]~35_combout ),
	.cout(\sReadCount[1]~36 ));
defparam \sReadCount[1]~35 .lut_mask = 16'h5A5F;
defparam \sReadCount[1]~35 .sum_lutc_input = "cin";

dffeas \sReadCount[1] (
	.clk(Clk),
	.d(\sReadCount[1]~35_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReadCount[0]~34_combout ),
	.q(\sReadCount[1]~q ),
	.prn(vcc));
defparam \sReadCount[1] .is_wysiwyg = "true";
defparam \sReadCount[1] .power_up = "low";

dffeas \sRegByteEnable[1] (
	.clk(Clk),
	.d(d_writedata_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sRegByteEnable[0]~2_combout ),
	.q(\sRegByteEnable[1]~q ),
	.prn(vcc));
defparam \sRegByteEnable[1] .is_wysiwyg = "true";
defparam \sRegByteEnable[1] .power_up = "low";

dffeas \sReg[1] (
	.clk(Clk),
	.d(d_writedata_1),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReg[0]~0_combout ),
	.q(\sReg[1]~q ),
	.prn(vcc));
defparam \sReg[1] .is_wysiwyg = "true";
defparam \sReg[1] .power_up = "low";

cycloneive_lcell_comb \ReadData[1]~2 (
	.dataa(W_alu_result_3),
	.datab(\sRegByteEnable[1]~q ),
	.datac(W_alu_result_2),
	.datad(\sReg[1]~q ),
	.cin(gnd),
	.combout(\ReadData[1]~2_combout ),
	.cout());
defparam \ReadData[1]~2 .lut_mask = 16'hFFDE;
defparam \ReadData[1]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sReadCountPipelined[1]~35 (
	.dataa(\sReadCountPipelined[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCountPipelined[0]~34 ),
	.combout(\sReadCountPipelined[1]~35_combout ),
	.cout(\sReadCountPipelined[1]~36 ));
defparam \sReadCountPipelined[1]~35 .lut_mask = 16'h5A5F;
defparam \sReadCountPipelined[1]~35 .sum_lutc_input = "cin";

dffeas \sReadCountPipelined[1] (
	.clk(Clk),
	.d(\sReadCountPipelined[1]~35_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sReadCountPipelined_0),
	.q(\sReadCountPipelined[1]~q ),
	.prn(vcc));
defparam \sReadCountPipelined[1] .is_wysiwyg = "true";
defparam \sReadCountPipelined[1] .power_up = "low";

dffeas \sRegByteEnable[2] (
	.clk(Clk),
	.d(d_writedata_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sRegByteEnable[0]~2_combout ),
	.q(\sRegByteEnable[2]~q ),
	.prn(vcc));
defparam \sRegByteEnable[2] .is_wysiwyg = "true";
defparam \sRegByteEnable[2] .power_up = "low";

cycloneive_lcell_comb \sReadCount[2]~37 (
	.dataa(\sReadCount[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCount[1]~36 ),
	.combout(\sReadCount[2]~37_combout ),
	.cout(\sReadCount[2]~38 ));
defparam \sReadCount[2]~37 .lut_mask = 16'h5AAF;
defparam \sReadCount[2]~37 .sum_lutc_input = "cin";

dffeas \sReadCount[2] (
	.clk(Clk),
	.d(\sReadCount[2]~37_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReadCount[0]~34_combout ),
	.q(\sReadCount[2]~q ),
	.prn(vcc));
defparam \sReadCount[2] .is_wysiwyg = "true";
defparam \sReadCount[2] .power_up = "low";

dffeas \sReg[2] (
	.clk(Clk),
	.d(d_writedata_2),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReg[0]~0_combout ),
	.q(\sReg[2]~q ),
	.prn(vcc));
defparam \sReg[2] .is_wysiwyg = "true";
defparam \sReg[2] .power_up = "low";

cycloneive_lcell_comb \ReadData[2]~4 (
	.dataa(W_alu_result_2),
	.datab(\sReadCount[2]~q ),
	.datac(W_alu_result_3),
	.datad(\sReg[2]~q ),
	.cin(gnd),
	.combout(\ReadData[2]~4_combout ),
	.cout());
defparam \ReadData[2]~4 .lut_mask = 16'hFFDE;
defparam \ReadData[2]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sReadCountPipelined[2]~37 (
	.dataa(\sReadCountPipelined[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCountPipelined[1]~36 ),
	.combout(\sReadCountPipelined[2]~37_combout ),
	.cout(\sReadCountPipelined[2]~38 ));
defparam \sReadCountPipelined[2]~37 .lut_mask = 16'h5AAF;
defparam \sReadCountPipelined[2]~37 .sum_lutc_input = "cin";

dffeas \sReadCountPipelined[2] (
	.clk(Clk),
	.d(\sReadCountPipelined[2]~37_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sReadCountPipelined_0),
	.q(\sReadCountPipelined[2]~q ),
	.prn(vcc));
defparam \sReadCountPipelined[2] .is_wysiwyg = "true";
defparam \sReadCountPipelined[2] .power_up = "low";

cycloneive_lcell_comb \sReadCount[3]~39 (
	.dataa(\sReadCount[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCount[2]~38 ),
	.combout(\sReadCount[3]~39_combout ),
	.cout(\sReadCount[3]~40 ));
defparam \sReadCount[3]~39 .lut_mask = 16'h5A5F;
defparam \sReadCount[3]~39 .sum_lutc_input = "cin";

dffeas \sReadCount[3] (
	.clk(Clk),
	.d(\sReadCount[3]~39_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReadCount[0]~34_combout ),
	.q(\sReadCount[3]~q ),
	.prn(vcc));
defparam \sReadCount[3] .is_wysiwyg = "true";
defparam \sReadCount[3] .power_up = "low";

dffeas \sRegByteEnable[3] (
	.clk(Clk),
	.d(d_writedata_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sRegByteEnable[0]~2_combout ),
	.q(\sRegByteEnable[3]~q ),
	.prn(vcc));
defparam \sRegByteEnable[3] .is_wysiwyg = "true";
defparam \sRegByteEnable[3] .power_up = "low";

dffeas \sReg[3] (
	.clk(Clk),
	.d(d_writedata_3),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReg[0]~0_combout ),
	.q(\sReg[3]~q ),
	.prn(vcc));
defparam \sReg[3] .is_wysiwyg = "true";
defparam \sReg[3] .power_up = "low";

cycloneive_lcell_comb \ReadData[3]~6 (
	.dataa(W_alu_result_3),
	.datab(\sRegByteEnable[3]~q ),
	.datac(W_alu_result_2),
	.datad(\sReg[3]~q ),
	.cin(gnd),
	.combout(\ReadData[3]~6_combout ),
	.cout());
defparam \ReadData[3]~6 .lut_mask = 16'hFFDE;
defparam \ReadData[3]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sReadCountPipelined[3]~39 (
	.dataa(\sReadCountPipelined[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCountPipelined[2]~38 ),
	.combout(\sReadCountPipelined[3]~39_combout ),
	.cout(\sReadCountPipelined[3]~40 ));
defparam \sReadCountPipelined[3]~39 .lut_mask = 16'h5A5F;
defparam \sReadCountPipelined[3]~39 .sum_lutc_input = "cin";

dffeas \sReadCountPipelined[3] (
	.clk(Clk),
	.d(\sReadCountPipelined[3]~39_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sReadCountPipelined_0),
	.q(\sReadCountPipelined[3]~q ),
	.prn(vcc));
defparam \sReadCountPipelined[3] .is_wysiwyg = "true";
defparam \sReadCountPipelined[3] .power_up = "low";

dffeas \sRegByteEnable[4] (
	.clk(Clk),
	.d(d_writedata_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sRegByteEnable[0]~2_combout ),
	.q(\sRegByteEnable[4]~q ),
	.prn(vcc));
defparam \sRegByteEnable[4] .is_wysiwyg = "true";
defparam \sRegByteEnable[4] .power_up = "low";

cycloneive_lcell_comb \sReadCount[4]~41 (
	.dataa(\sReadCount[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCount[3]~40 ),
	.combout(\sReadCount[4]~41_combout ),
	.cout(\sReadCount[4]~42 ));
defparam \sReadCount[4]~41 .lut_mask = 16'h5AAF;
defparam \sReadCount[4]~41 .sum_lutc_input = "cin";

dffeas \sReadCount[4] (
	.clk(Clk),
	.d(\sReadCount[4]~41_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReadCount[0]~34_combout ),
	.q(\sReadCount[4]~q ),
	.prn(vcc));
defparam \sReadCount[4] .is_wysiwyg = "true";
defparam \sReadCount[4] .power_up = "low";

dffeas \sReg[4] (
	.clk(Clk),
	.d(d_writedata_4),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReg[0]~0_combout ),
	.q(\sReg[4]~q ),
	.prn(vcc));
defparam \sReg[4] .is_wysiwyg = "true";
defparam \sReg[4] .power_up = "low";

cycloneive_lcell_comb \ReadData[4]~8 (
	.dataa(W_alu_result_2),
	.datab(\sReadCount[4]~q ),
	.datac(W_alu_result_3),
	.datad(\sReg[4]~q ),
	.cin(gnd),
	.combout(\ReadData[4]~8_combout ),
	.cout());
defparam \ReadData[4]~8 .lut_mask = 16'hFFDE;
defparam \ReadData[4]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sReadCountPipelined[4]~41 (
	.dataa(\sReadCountPipelined[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCountPipelined[3]~40 ),
	.combout(\sReadCountPipelined[4]~41_combout ),
	.cout(\sReadCountPipelined[4]~42 ));
defparam \sReadCountPipelined[4]~41 .lut_mask = 16'h5AAF;
defparam \sReadCountPipelined[4]~41 .sum_lutc_input = "cin";

dffeas \sReadCountPipelined[4] (
	.clk(Clk),
	.d(\sReadCountPipelined[4]~41_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sReadCountPipelined_0),
	.q(\sReadCountPipelined[4]~q ),
	.prn(vcc));
defparam \sReadCountPipelined[4] .is_wysiwyg = "true";
defparam \sReadCountPipelined[4] .power_up = "low";

cycloneive_lcell_comb \sReadCount[5]~43 (
	.dataa(\sReadCount[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCount[4]~42 ),
	.combout(\sReadCount[5]~43_combout ),
	.cout(\sReadCount[5]~44 ));
defparam \sReadCount[5]~43 .lut_mask = 16'h5A5F;
defparam \sReadCount[5]~43 .sum_lutc_input = "cin";

dffeas \sReadCount[5] (
	.clk(Clk),
	.d(\sReadCount[5]~43_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReadCount[0]~34_combout ),
	.q(\sReadCount[5]~q ),
	.prn(vcc));
defparam \sReadCount[5] .is_wysiwyg = "true";
defparam \sReadCount[5] .power_up = "low";

dffeas \sRegByteEnable[5] (
	.clk(Clk),
	.d(d_writedata_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sRegByteEnable[0]~2_combout ),
	.q(\sRegByteEnable[5]~q ),
	.prn(vcc));
defparam \sRegByteEnable[5] .is_wysiwyg = "true";
defparam \sRegByteEnable[5] .power_up = "low";

dffeas \sReg[5] (
	.clk(Clk),
	.d(d_writedata_5),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReg[0]~0_combout ),
	.q(\sReg[5]~q ),
	.prn(vcc));
defparam \sReg[5] .is_wysiwyg = "true";
defparam \sReg[5] .power_up = "low";

cycloneive_lcell_comb \ReadData[5]~10 (
	.dataa(W_alu_result_3),
	.datab(\sRegByteEnable[5]~q ),
	.datac(W_alu_result_2),
	.datad(\sReg[5]~q ),
	.cin(gnd),
	.combout(\ReadData[5]~10_combout ),
	.cout());
defparam \ReadData[5]~10 .lut_mask = 16'hFFDE;
defparam \ReadData[5]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sReadCountPipelined[5]~43 (
	.dataa(\sReadCountPipelined[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCountPipelined[4]~42 ),
	.combout(\sReadCountPipelined[5]~43_combout ),
	.cout(\sReadCountPipelined[5]~44 ));
defparam \sReadCountPipelined[5]~43 .lut_mask = 16'h5A5F;
defparam \sReadCountPipelined[5]~43 .sum_lutc_input = "cin";

dffeas \sReadCountPipelined[5] (
	.clk(Clk),
	.d(\sReadCountPipelined[5]~43_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sReadCountPipelined_0),
	.q(\sReadCountPipelined[5]~q ),
	.prn(vcc));
defparam \sReadCountPipelined[5] .is_wysiwyg = "true";
defparam \sReadCountPipelined[5] .power_up = "low";

dffeas \sRegByteEnable[6] (
	.clk(Clk),
	.d(d_writedata_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sRegByteEnable[0]~2_combout ),
	.q(\sRegByteEnable[6]~q ),
	.prn(vcc));
defparam \sRegByteEnable[6] .is_wysiwyg = "true";
defparam \sRegByteEnable[6] .power_up = "low";

cycloneive_lcell_comb \sReadCount[6]~45 (
	.dataa(\sReadCount[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCount[5]~44 ),
	.combout(\sReadCount[6]~45_combout ),
	.cout(\sReadCount[6]~46 ));
defparam \sReadCount[6]~45 .lut_mask = 16'h5AAF;
defparam \sReadCount[6]~45 .sum_lutc_input = "cin";

dffeas \sReadCount[6] (
	.clk(Clk),
	.d(\sReadCount[6]~45_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReadCount[0]~34_combout ),
	.q(\sReadCount[6]~q ),
	.prn(vcc));
defparam \sReadCount[6] .is_wysiwyg = "true";
defparam \sReadCount[6] .power_up = "low";

dffeas \sReg[6] (
	.clk(Clk),
	.d(d_writedata_6),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReg[0]~0_combout ),
	.q(\sReg[6]~q ),
	.prn(vcc));
defparam \sReg[6] .is_wysiwyg = "true";
defparam \sReg[6] .power_up = "low";

cycloneive_lcell_comb \ReadData[6]~12 (
	.dataa(W_alu_result_2),
	.datab(\sReadCount[6]~q ),
	.datac(W_alu_result_3),
	.datad(\sReg[6]~q ),
	.cin(gnd),
	.combout(\ReadData[6]~12_combout ),
	.cout());
defparam \ReadData[6]~12 .lut_mask = 16'hFFDE;
defparam \ReadData[6]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sReadCountPipelined[6]~45 (
	.dataa(\sReadCountPipelined[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCountPipelined[5]~44 ),
	.combout(\sReadCountPipelined[6]~45_combout ),
	.cout(\sReadCountPipelined[6]~46 ));
defparam \sReadCountPipelined[6]~45 .lut_mask = 16'h5AAF;
defparam \sReadCountPipelined[6]~45 .sum_lutc_input = "cin";

dffeas \sReadCountPipelined[6] (
	.clk(Clk),
	.d(\sReadCountPipelined[6]~45_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sReadCountPipelined_0),
	.q(\sReadCountPipelined[6]~q ),
	.prn(vcc));
defparam \sReadCountPipelined[6] .is_wysiwyg = "true";
defparam \sReadCountPipelined[6] .power_up = "low";

cycloneive_lcell_comb \sReadCount[7]~47 (
	.dataa(\sReadCount[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCount[6]~46 ),
	.combout(\sReadCount[7]~47_combout ),
	.cout(\sReadCount[7]~48 ));
defparam \sReadCount[7]~47 .lut_mask = 16'h5A5F;
defparam \sReadCount[7]~47 .sum_lutc_input = "cin";

dffeas \sReadCount[7] (
	.clk(Clk),
	.d(\sReadCount[7]~47_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReadCount[0]~34_combout ),
	.q(\sReadCount[7]~q ),
	.prn(vcc));
defparam \sReadCount[7] .is_wysiwyg = "true";
defparam \sReadCount[7] .power_up = "low";

dffeas \sRegByteEnable[7] (
	.clk(Clk),
	.d(d_writedata_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sRegByteEnable[0]~2_combout ),
	.q(\sRegByteEnable[7]~q ),
	.prn(vcc));
defparam \sRegByteEnable[7] .is_wysiwyg = "true";
defparam \sRegByteEnable[7] .power_up = "low";

dffeas \sReg[7] (
	.clk(Clk),
	.d(d_writedata_7),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReg[0]~0_combout ),
	.q(\sReg[7]~q ),
	.prn(vcc));
defparam \sReg[7] .is_wysiwyg = "true";
defparam \sReg[7] .power_up = "low";

cycloneive_lcell_comb \ReadData[7]~14 (
	.dataa(W_alu_result_3),
	.datab(\sRegByteEnable[7]~q ),
	.datac(W_alu_result_2),
	.datad(\sReg[7]~q ),
	.cin(gnd),
	.combout(\ReadData[7]~14_combout ),
	.cout());
defparam \ReadData[7]~14 .lut_mask = 16'hFFDE;
defparam \ReadData[7]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sReadCountPipelined[7]~47 (
	.dataa(\sReadCountPipelined[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCountPipelined[6]~46 ),
	.combout(\sReadCountPipelined[7]~47_combout ),
	.cout(\sReadCountPipelined[7]~48 ));
defparam \sReadCountPipelined[7]~47 .lut_mask = 16'h5A5F;
defparam \sReadCountPipelined[7]~47 .sum_lutc_input = "cin";

dffeas \sReadCountPipelined[7] (
	.clk(Clk),
	.d(\sReadCountPipelined[7]~47_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sReadCountPipelined_0),
	.q(\sReadCountPipelined[7]~q ),
	.prn(vcc));
defparam \sReadCountPipelined[7] .is_wysiwyg = "true";
defparam \sReadCountPipelined[7] .power_up = "low";

cycloneive_lcell_comb \sRegByteEnable[8]~3 (
	.dataa(d_byteenable_1),
	.datab(\sRegByteEnable[24]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sRegByteEnable[8]~3_combout ),
	.cout());
defparam \sRegByteEnable[8]~3 .lut_mask = 16'hEEEE;
defparam \sRegByteEnable[8]~3 .sum_lutc_input = "datac";

dffeas \sRegByteEnable[8] (
	.clk(Clk),
	.d(d_writedata_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sRegByteEnable[8]~3_combout ),
	.q(\sRegByteEnable[8]~q ),
	.prn(vcc));
defparam \sRegByteEnable[8] .is_wysiwyg = "true";
defparam \sRegByteEnable[8] .power_up = "low";

cycloneive_lcell_comb \sReadCount[8]~49 (
	.dataa(\sReadCount[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCount[7]~48 ),
	.combout(\sReadCount[8]~49_combout ),
	.cout(\sReadCount[8]~50 ));
defparam \sReadCount[8]~49 .lut_mask = 16'h5AAF;
defparam \sReadCount[8]~49 .sum_lutc_input = "cin";

dffeas \sReadCount[8] (
	.clk(Clk),
	.d(\sReadCount[8]~49_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReadCount[0]~34_combout ),
	.q(\sReadCount[8]~q ),
	.prn(vcc));
defparam \sReadCount[8] .is_wysiwyg = "true";
defparam \sReadCount[8] .power_up = "low";

dffeas \sReg[8] (
	.clk(Clk),
	.d(d_writedata_8),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReg[0]~0_combout ),
	.q(\sReg[8]~q ),
	.prn(vcc));
defparam \sReg[8] .is_wysiwyg = "true";
defparam \sReg[8] .power_up = "low";

cycloneive_lcell_comb \ReadData[8]~16 (
	.dataa(W_alu_result_2),
	.datab(\sReadCount[8]~q ),
	.datac(W_alu_result_3),
	.datad(\sReg[8]~q ),
	.cin(gnd),
	.combout(\ReadData[8]~16_combout ),
	.cout());
defparam \ReadData[8]~16 .lut_mask = 16'hFFDE;
defparam \ReadData[8]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sReadCountPipelined[8]~49 (
	.dataa(\sReadCountPipelined[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCountPipelined[7]~48 ),
	.combout(\sReadCountPipelined[8]~49_combout ),
	.cout(\sReadCountPipelined[8]~50 ));
defparam \sReadCountPipelined[8]~49 .lut_mask = 16'h5AAF;
defparam \sReadCountPipelined[8]~49 .sum_lutc_input = "cin";

dffeas \sReadCountPipelined[8] (
	.clk(Clk),
	.d(\sReadCountPipelined[8]~49_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sReadCountPipelined_0),
	.q(\sReadCountPipelined[8]~q ),
	.prn(vcc));
defparam \sReadCountPipelined[8] .is_wysiwyg = "true";
defparam \sReadCountPipelined[8] .power_up = "low";

dffeas \sRegByteEnable[12] (
	.clk(Clk),
	.d(d_writedata_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sRegByteEnable[8]~3_combout ),
	.q(\sRegByteEnable[12]~q ),
	.prn(vcc));
defparam \sRegByteEnable[12] .is_wysiwyg = "true";
defparam \sRegByteEnable[12] .power_up = "low";

cycloneive_lcell_comb \sReadCount[9]~51 (
	.dataa(\sReadCount[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCount[8]~50 ),
	.combout(\sReadCount[9]~51_combout ),
	.cout(\sReadCount[9]~52 ));
defparam \sReadCount[9]~51 .lut_mask = 16'h5A5F;
defparam \sReadCount[9]~51 .sum_lutc_input = "cin";

dffeas \sReadCount[9] (
	.clk(Clk),
	.d(\sReadCount[9]~51_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReadCount[0]~34_combout ),
	.q(\sReadCount[9]~q ),
	.prn(vcc));
defparam \sReadCount[9] .is_wysiwyg = "true";
defparam \sReadCount[9] .power_up = "low";

cycloneive_lcell_comb \sReadCount[10]~53 (
	.dataa(\sReadCount[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCount[9]~52 ),
	.combout(\sReadCount[10]~53_combout ),
	.cout(\sReadCount[10]~54 ));
defparam \sReadCount[10]~53 .lut_mask = 16'h5AAF;
defparam \sReadCount[10]~53 .sum_lutc_input = "cin";

dffeas \sReadCount[10] (
	.clk(Clk),
	.d(\sReadCount[10]~53_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReadCount[0]~34_combout ),
	.q(\sReadCount[10]~q ),
	.prn(vcc));
defparam \sReadCount[10] .is_wysiwyg = "true";
defparam \sReadCount[10] .power_up = "low";

cycloneive_lcell_comb \sReadCount[11]~55 (
	.dataa(\sReadCount[11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCount[10]~54 ),
	.combout(\sReadCount[11]~55_combout ),
	.cout(\sReadCount[11]~56 ));
defparam \sReadCount[11]~55 .lut_mask = 16'h5A5F;
defparam \sReadCount[11]~55 .sum_lutc_input = "cin";

dffeas \sReadCount[11] (
	.clk(Clk),
	.d(\sReadCount[11]~55_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReadCount[0]~34_combout ),
	.q(\sReadCount[11]~q ),
	.prn(vcc));
defparam \sReadCount[11] .is_wysiwyg = "true";
defparam \sReadCount[11] .power_up = "low";

cycloneive_lcell_comb \sReadCount[12]~57 (
	.dataa(\sReadCount[12]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCount[11]~56 ),
	.combout(\sReadCount[12]~57_combout ),
	.cout(\sReadCount[12]~58 ));
defparam \sReadCount[12]~57 .lut_mask = 16'h5AAF;
defparam \sReadCount[12]~57 .sum_lutc_input = "cin";

dffeas \sReadCount[12] (
	.clk(Clk),
	.d(\sReadCount[12]~57_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReadCount[0]~34_combout ),
	.q(\sReadCount[12]~q ),
	.prn(vcc));
defparam \sReadCount[12] .is_wysiwyg = "true";
defparam \sReadCount[12] .power_up = "low";

dffeas \sReg[12] (
	.clk(Clk),
	.d(d_writedata_12),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReg[0]~0_combout ),
	.q(\sReg[12]~q ),
	.prn(vcc));
defparam \sReg[12] .is_wysiwyg = "true";
defparam \sReg[12] .power_up = "low";

cycloneive_lcell_comb \ReadData[12]~18 (
	.dataa(W_alu_result_2),
	.datab(\sReadCount[12]~q ),
	.datac(W_alu_result_3),
	.datad(\sReg[12]~q ),
	.cin(gnd),
	.combout(\ReadData[12]~18_combout ),
	.cout());
defparam \ReadData[12]~18 .lut_mask = 16'hFFDE;
defparam \ReadData[12]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sReadCountPipelined[9]~51 (
	.dataa(\sReadCountPipelined[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCountPipelined[8]~50 ),
	.combout(\sReadCountPipelined[9]~51_combout ),
	.cout(\sReadCountPipelined[9]~52 ));
defparam \sReadCountPipelined[9]~51 .lut_mask = 16'h5A5F;
defparam \sReadCountPipelined[9]~51 .sum_lutc_input = "cin";

dffeas \sReadCountPipelined[9] (
	.clk(Clk),
	.d(\sReadCountPipelined[9]~51_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sReadCountPipelined_0),
	.q(\sReadCountPipelined[9]~q ),
	.prn(vcc));
defparam \sReadCountPipelined[9] .is_wysiwyg = "true";
defparam \sReadCountPipelined[9] .power_up = "low";

cycloneive_lcell_comb \sReadCountPipelined[10]~53 (
	.dataa(\sReadCountPipelined[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCountPipelined[9]~52 ),
	.combout(\sReadCountPipelined[10]~53_combout ),
	.cout(\sReadCountPipelined[10]~54 ));
defparam \sReadCountPipelined[10]~53 .lut_mask = 16'h5AAF;
defparam \sReadCountPipelined[10]~53 .sum_lutc_input = "cin";

dffeas \sReadCountPipelined[10] (
	.clk(Clk),
	.d(\sReadCountPipelined[10]~53_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sReadCountPipelined_0),
	.q(\sReadCountPipelined[10]~q ),
	.prn(vcc));
defparam \sReadCountPipelined[10] .is_wysiwyg = "true";
defparam \sReadCountPipelined[10] .power_up = "low";

cycloneive_lcell_comb \sReadCountPipelined[11]~55 (
	.dataa(\sReadCountPipelined[11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCountPipelined[10]~54 ),
	.combout(\sReadCountPipelined[11]~55_combout ),
	.cout(\sReadCountPipelined[11]~56 ));
defparam \sReadCountPipelined[11]~55 .lut_mask = 16'h5A5F;
defparam \sReadCountPipelined[11]~55 .sum_lutc_input = "cin";

dffeas \sReadCountPipelined[11] (
	.clk(Clk),
	.d(\sReadCountPipelined[11]~55_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sReadCountPipelined_0),
	.q(\sReadCountPipelined[11]~q ),
	.prn(vcc));
defparam \sReadCountPipelined[11] .is_wysiwyg = "true";
defparam \sReadCountPipelined[11] .power_up = "low";

cycloneive_lcell_comb \sReadCountPipelined[12]~57 (
	.dataa(\sReadCountPipelined[12]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCountPipelined[11]~56 ),
	.combout(\sReadCountPipelined[12]~57_combout ),
	.cout(\sReadCountPipelined[12]~58 ));
defparam \sReadCountPipelined[12]~57 .lut_mask = 16'h5AAF;
defparam \sReadCountPipelined[12]~57 .sum_lutc_input = "cin";

dffeas \sReadCountPipelined[12] (
	.clk(Clk),
	.d(\sReadCountPipelined[12]~57_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sReadCountPipelined_0),
	.q(\sReadCountPipelined[12]~q ),
	.prn(vcc));
defparam \sReadCountPipelined[12] .is_wysiwyg = "true";
defparam \sReadCountPipelined[12] .power_up = "low";

dffeas \sRegByteEnable[11] (
	.clk(Clk),
	.d(d_writedata_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sRegByteEnable[8]~3_combout ),
	.q(\sRegByteEnable[11]~q ),
	.prn(vcc));
defparam \sRegByteEnable[11] .is_wysiwyg = "true";
defparam \sRegByteEnable[11] .power_up = "low";

dffeas \sReg[11] (
	.clk(Clk),
	.d(d_writedata_11),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReg[0]~0_combout ),
	.q(\sReg[11]~q ),
	.prn(vcc));
defparam \sReg[11] .is_wysiwyg = "true";
defparam \sReg[11] .power_up = "low";

cycloneive_lcell_comb \ReadData[11]~20 (
	.dataa(W_alu_result_3),
	.datab(\sRegByteEnable[11]~q ),
	.datac(W_alu_result_2),
	.datad(\sReg[11]~q ),
	.cin(gnd),
	.combout(\ReadData[11]~20_combout ),
	.cout());
defparam \ReadData[11]~20 .lut_mask = 16'hFFDE;
defparam \ReadData[11]~20 .sum_lutc_input = "datac";

dffeas \sRegByteEnable[10] (
	.clk(Clk),
	.d(d_writedata_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sRegByteEnable[8]~3_combout ),
	.q(\sRegByteEnable[10]~q ),
	.prn(vcc));
defparam \sRegByteEnable[10] .is_wysiwyg = "true";
defparam \sRegByteEnable[10] .power_up = "low";

dffeas \sReg[10] (
	.clk(Clk),
	.d(d_writedata_10),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReg[0]~0_combout ),
	.q(\sReg[10]~q ),
	.prn(vcc));
defparam \sReg[10] .is_wysiwyg = "true";
defparam \sReg[10] .power_up = "low";

cycloneive_lcell_comb \ReadData[10]~22 (
	.dataa(W_alu_result_2),
	.datab(\sReadCount[10]~q ),
	.datac(W_alu_result_3),
	.datad(\sReg[10]~q ),
	.cin(gnd),
	.combout(\ReadData[10]~22_combout ),
	.cout());
defparam \ReadData[10]~22 .lut_mask = 16'hFFDE;
defparam \ReadData[10]~22 .sum_lutc_input = "datac";

dffeas \sRegByteEnable[9] (
	.clk(Clk),
	.d(d_writedata_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sRegByteEnable[8]~3_combout ),
	.q(\sRegByteEnable[9]~q ),
	.prn(vcc));
defparam \sRegByteEnable[9] .is_wysiwyg = "true";
defparam \sRegByteEnable[9] .power_up = "low";

dffeas \sReg[9] (
	.clk(Clk),
	.d(d_writedata_9),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReg[0]~0_combout ),
	.q(\sReg[9]~q ),
	.prn(vcc));
defparam \sReg[9] .is_wysiwyg = "true";
defparam \sReg[9] .power_up = "low";

cycloneive_lcell_comb \ReadData[9]~24 (
	.dataa(W_alu_result_3),
	.datab(\sRegByteEnable[9]~q ),
	.datac(W_alu_result_2),
	.datad(\sReg[9]~q ),
	.cin(gnd),
	.combout(\ReadData[9]~24_combout ),
	.cout());
defparam \ReadData[9]~24 .lut_mask = 16'hFFDE;
defparam \ReadData[9]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sReadCount[13]~59 (
	.dataa(\sReadCount[13]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCount[12]~58 ),
	.combout(\sReadCount[13]~59_combout ),
	.cout(\sReadCount[13]~60 ));
defparam \sReadCount[13]~59 .lut_mask = 16'h5A5F;
defparam \sReadCount[13]~59 .sum_lutc_input = "cin";

dffeas \sReadCount[13] (
	.clk(Clk),
	.d(\sReadCount[13]~59_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReadCount[0]~34_combout ),
	.q(\sReadCount[13]~q ),
	.prn(vcc));
defparam \sReadCount[13] .is_wysiwyg = "true";
defparam \sReadCount[13] .power_up = "low";

cycloneive_lcell_comb \sReadCount[14]~61 (
	.dataa(\sReadCount[14]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCount[13]~60 ),
	.combout(\sReadCount[14]~61_combout ),
	.cout(\sReadCount[14]~62 ));
defparam \sReadCount[14]~61 .lut_mask = 16'h5AAF;
defparam \sReadCount[14]~61 .sum_lutc_input = "cin";

dffeas \sReadCount[14] (
	.clk(Clk),
	.d(\sReadCount[14]~61_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReadCount[0]~34_combout ),
	.q(\sReadCount[14]~q ),
	.prn(vcc));
defparam \sReadCount[14] .is_wysiwyg = "true";
defparam \sReadCount[14] .power_up = "low";

cycloneive_lcell_comb \sReadCount[15]~63 (
	.dataa(\sReadCount[15]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCount[14]~62 ),
	.combout(\sReadCount[15]~63_combout ),
	.cout(\sReadCount[15]~64 ));
defparam \sReadCount[15]~63 .lut_mask = 16'h5A5F;
defparam \sReadCount[15]~63 .sum_lutc_input = "cin";

dffeas \sReadCount[15] (
	.clk(Clk),
	.d(\sReadCount[15]~63_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReadCount[0]~34_combout ),
	.q(\sReadCount[15]~q ),
	.prn(vcc));
defparam \sReadCount[15] .is_wysiwyg = "true";
defparam \sReadCount[15] .power_up = "low";

dffeas \sRegByteEnable[15] (
	.clk(Clk),
	.d(d_writedata_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sRegByteEnable[8]~3_combout ),
	.q(\sRegByteEnable[15]~q ),
	.prn(vcc));
defparam \sRegByteEnable[15] .is_wysiwyg = "true";
defparam \sRegByteEnable[15] .power_up = "low";

dffeas \sReg[15] (
	.clk(Clk),
	.d(d_writedata_15),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReg[0]~0_combout ),
	.q(\sReg[15]~q ),
	.prn(vcc));
defparam \sReg[15] .is_wysiwyg = "true";
defparam \sReg[15] .power_up = "low";

cycloneive_lcell_comb \ReadData[15]~26 (
	.dataa(W_alu_result_3),
	.datab(\sRegByteEnable[15]~q ),
	.datac(W_alu_result_2),
	.datad(\sReg[15]~q ),
	.cin(gnd),
	.combout(\ReadData[15]~26_combout ),
	.cout());
defparam \ReadData[15]~26 .lut_mask = 16'hFFDE;
defparam \ReadData[15]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sReadCountPipelined[13]~59 (
	.dataa(\sReadCountPipelined[13]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCountPipelined[12]~58 ),
	.combout(\sReadCountPipelined[13]~59_combout ),
	.cout(\sReadCountPipelined[13]~60 ));
defparam \sReadCountPipelined[13]~59 .lut_mask = 16'h5A5F;
defparam \sReadCountPipelined[13]~59 .sum_lutc_input = "cin";

dffeas \sReadCountPipelined[13] (
	.clk(Clk),
	.d(\sReadCountPipelined[13]~59_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sReadCountPipelined_0),
	.q(\sReadCountPipelined[13]~q ),
	.prn(vcc));
defparam \sReadCountPipelined[13] .is_wysiwyg = "true";
defparam \sReadCountPipelined[13] .power_up = "low";

cycloneive_lcell_comb \sReadCountPipelined[14]~61 (
	.dataa(\sReadCountPipelined[14]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCountPipelined[13]~60 ),
	.combout(\sReadCountPipelined[14]~61_combout ),
	.cout(\sReadCountPipelined[14]~62 ));
defparam \sReadCountPipelined[14]~61 .lut_mask = 16'h5AAF;
defparam \sReadCountPipelined[14]~61 .sum_lutc_input = "cin";

dffeas \sReadCountPipelined[14] (
	.clk(Clk),
	.d(\sReadCountPipelined[14]~61_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sReadCountPipelined_0),
	.q(\sReadCountPipelined[14]~q ),
	.prn(vcc));
defparam \sReadCountPipelined[14] .is_wysiwyg = "true";
defparam \sReadCountPipelined[14] .power_up = "low";

cycloneive_lcell_comb \sReadCountPipelined[15]~63 (
	.dataa(\sReadCountPipelined[15]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCountPipelined[14]~62 ),
	.combout(\sReadCountPipelined[15]~63_combout ),
	.cout(\sReadCountPipelined[15]~64 ));
defparam \sReadCountPipelined[15]~63 .lut_mask = 16'h5A5F;
defparam \sReadCountPipelined[15]~63 .sum_lutc_input = "cin";

dffeas \sReadCountPipelined[15] (
	.clk(Clk),
	.d(\sReadCountPipelined[15]~63_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sReadCountPipelined_0),
	.q(\sReadCountPipelined[15]~q ),
	.prn(vcc));
defparam \sReadCountPipelined[15] .is_wysiwyg = "true";
defparam \sReadCountPipelined[15] .power_up = "low";

dffeas \sRegByteEnable[14] (
	.clk(Clk),
	.d(d_writedata_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sRegByteEnable[8]~3_combout ),
	.q(\sRegByteEnable[14]~q ),
	.prn(vcc));
defparam \sRegByteEnable[14] .is_wysiwyg = "true";
defparam \sRegByteEnable[14] .power_up = "low";

dffeas \sReg[14] (
	.clk(Clk),
	.d(d_writedata_14),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReg[0]~0_combout ),
	.q(\sReg[14]~q ),
	.prn(vcc));
defparam \sReg[14] .is_wysiwyg = "true";
defparam \sReg[14] .power_up = "low";

cycloneive_lcell_comb \ReadData[14]~28 (
	.dataa(W_alu_result_2),
	.datab(\sReadCount[14]~q ),
	.datac(W_alu_result_3),
	.datad(\sReg[14]~q ),
	.cin(gnd),
	.combout(\ReadData[14]~28_combout ),
	.cout());
defparam \ReadData[14]~28 .lut_mask = 16'hFFDE;
defparam \ReadData[14]~28 .sum_lutc_input = "datac";

dffeas \sRegByteEnable[13] (
	.clk(Clk),
	.d(d_writedata_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sRegByteEnable[8]~3_combout ),
	.q(\sRegByteEnable[13]~q ),
	.prn(vcc));
defparam \sRegByteEnable[13] .is_wysiwyg = "true";
defparam \sRegByteEnable[13] .power_up = "low";

dffeas \sReg[13] (
	.clk(Clk),
	.d(d_writedata_13),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReg[0]~0_combout ),
	.q(\sReg[13]~q ),
	.prn(vcc));
defparam \sReg[13] .is_wysiwyg = "true";
defparam \sReg[13] .power_up = "low";

cycloneive_lcell_comb \ReadData[13]~30 (
	.dataa(W_alu_result_3),
	.datab(\sRegByteEnable[13]~q ),
	.datac(W_alu_result_2),
	.datad(\sReg[13]~q ),
	.cin(gnd),
	.combout(\ReadData[13]~30_combout ),
	.cout());
defparam \ReadData[13]~30 .lut_mask = 16'hFFDE;
defparam \ReadData[13]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sRegByteEnable[16]~4 (
	.dataa(d_byteenable_2),
	.datab(\sRegByteEnable[24]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sRegByteEnable[16]~4_combout ),
	.cout());
defparam \sRegByteEnable[16]~4 .lut_mask = 16'hEEEE;
defparam \sRegByteEnable[16]~4 .sum_lutc_input = "datac";

dffeas \sRegByteEnable[16] (
	.clk(Clk),
	.d(d_writedata_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sRegByteEnable[16]~4_combout ),
	.q(\sRegByteEnable[16]~q ),
	.prn(vcc));
defparam \sRegByteEnable[16] .is_wysiwyg = "true";
defparam \sRegByteEnable[16] .power_up = "low";

cycloneive_lcell_comb \sReadCount[16]~65 (
	.dataa(\sReadCount[16]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCount[15]~64 ),
	.combout(\sReadCount[16]~65_combout ),
	.cout(\sReadCount[16]~66 ));
defparam \sReadCount[16]~65 .lut_mask = 16'h5AAF;
defparam \sReadCount[16]~65 .sum_lutc_input = "cin";

dffeas \sReadCount[16] (
	.clk(Clk),
	.d(\sReadCount[16]~65_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReadCount[0]~34_combout ),
	.q(\sReadCount[16]~q ),
	.prn(vcc));
defparam \sReadCount[16] .is_wysiwyg = "true";
defparam \sReadCount[16] .power_up = "low";

dffeas \sReg[16] (
	.clk(Clk),
	.d(d_writedata_16),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReg[0]~0_combout ),
	.q(\sReg[16]~q ),
	.prn(vcc));
defparam \sReg[16] .is_wysiwyg = "true";
defparam \sReg[16] .power_up = "low";

cycloneive_lcell_comb \ReadData[16]~32 (
	.dataa(W_alu_result_2),
	.datab(\sReadCount[16]~q ),
	.datac(W_alu_result_3),
	.datad(\sReg[16]~q ),
	.cin(gnd),
	.combout(\ReadData[16]~32_combout ),
	.cout());
defparam \ReadData[16]~32 .lut_mask = 16'hFFDE;
defparam \ReadData[16]~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sReadCountPipelined[16]~65 (
	.dataa(\sReadCountPipelined[16]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCountPipelined[15]~64 ),
	.combout(\sReadCountPipelined[16]~65_combout ),
	.cout(\sReadCountPipelined[16]~66 ));
defparam \sReadCountPipelined[16]~65 .lut_mask = 16'h5AAF;
defparam \sReadCountPipelined[16]~65 .sum_lutc_input = "cin";

dffeas \sReadCountPipelined[16] (
	.clk(Clk),
	.d(\sReadCountPipelined[16]~65_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sReadCountPipelined_0),
	.q(\sReadCountPipelined[16]~q ),
	.prn(vcc));
defparam \sReadCountPipelined[16] .is_wysiwyg = "true";
defparam \sReadCountPipelined[16] .power_up = "low";

dffeas \sRegByteEnable[20] (
	.clk(Clk),
	.d(d_writedata_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sRegByteEnable[16]~4_combout ),
	.q(\sRegByteEnable[20]~q ),
	.prn(vcc));
defparam \sRegByteEnable[20] .is_wysiwyg = "true";
defparam \sRegByteEnable[20] .power_up = "low";

cycloneive_lcell_comb \sReadCount[17]~67 (
	.dataa(\sReadCount[17]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCount[16]~66 ),
	.combout(\sReadCount[17]~67_combout ),
	.cout(\sReadCount[17]~68 ));
defparam \sReadCount[17]~67 .lut_mask = 16'h5A5F;
defparam \sReadCount[17]~67 .sum_lutc_input = "cin";

dffeas \sReadCount[17] (
	.clk(Clk),
	.d(\sReadCount[17]~67_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReadCount[0]~34_combout ),
	.q(\sReadCount[17]~q ),
	.prn(vcc));
defparam \sReadCount[17] .is_wysiwyg = "true";
defparam \sReadCount[17] .power_up = "low";

cycloneive_lcell_comb \sReadCount[18]~69 (
	.dataa(\sReadCount[18]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCount[17]~68 ),
	.combout(\sReadCount[18]~69_combout ),
	.cout(\sReadCount[18]~70 ));
defparam \sReadCount[18]~69 .lut_mask = 16'h5AAF;
defparam \sReadCount[18]~69 .sum_lutc_input = "cin";

dffeas \sReadCount[18] (
	.clk(Clk),
	.d(\sReadCount[18]~69_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReadCount[0]~34_combout ),
	.q(\sReadCount[18]~q ),
	.prn(vcc));
defparam \sReadCount[18] .is_wysiwyg = "true";
defparam \sReadCount[18] .power_up = "low";

cycloneive_lcell_comb \sReadCount[19]~71 (
	.dataa(\sReadCount[19]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCount[18]~70 ),
	.combout(\sReadCount[19]~71_combout ),
	.cout(\sReadCount[19]~72 ));
defparam \sReadCount[19]~71 .lut_mask = 16'h5A5F;
defparam \sReadCount[19]~71 .sum_lutc_input = "cin";

dffeas \sReadCount[19] (
	.clk(Clk),
	.d(\sReadCount[19]~71_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReadCount[0]~34_combout ),
	.q(\sReadCount[19]~q ),
	.prn(vcc));
defparam \sReadCount[19] .is_wysiwyg = "true";
defparam \sReadCount[19] .power_up = "low";

cycloneive_lcell_comb \sReadCount[20]~73 (
	.dataa(\sReadCount[20]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCount[19]~72 ),
	.combout(\sReadCount[20]~73_combout ),
	.cout(\sReadCount[20]~74 ));
defparam \sReadCount[20]~73 .lut_mask = 16'h5AAF;
defparam \sReadCount[20]~73 .sum_lutc_input = "cin";

dffeas \sReadCount[20] (
	.clk(Clk),
	.d(\sReadCount[20]~73_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReadCount[0]~34_combout ),
	.q(\sReadCount[20]~q ),
	.prn(vcc));
defparam \sReadCount[20] .is_wysiwyg = "true";
defparam \sReadCount[20] .power_up = "low";

dffeas \sReg[20] (
	.clk(Clk),
	.d(d_writedata_20),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReg[0]~0_combout ),
	.q(\sReg[20]~q ),
	.prn(vcc));
defparam \sReg[20] .is_wysiwyg = "true";
defparam \sReg[20] .power_up = "low";

cycloneive_lcell_comb \ReadData[20]~34 (
	.dataa(W_alu_result_2),
	.datab(\sReadCount[20]~q ),
	.datac(W_alu_result_3),
	.datad(\sReg[20]~q ),
	.cin(gnd),
	.combout(\ReadData[20]~34_combout ),
	.cout());
defparam \ReadData[20]~34 .lut_mask = 16'hFFDE;
defparam \ReadData[20]~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sReadCountPipelined[17]~67 (
	.dataa(\sReadCountPipelined[17]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCountPipelined[16]~66 ),
	.combout(\sReadCountPipelined[17]~67_combout ),
	.cout(\sReadCountPipelined[17]~68 ));
defparam \sReadCountPipelined[17]~67 .lut_mask = 16'h5A5F;
defparam \sReadCountPipelined[17]~67 .sum_lutc_input = "cin";

dffeas \sReadCountPipelined[17] (
	.clk(Clk),
	.d(\sReadCountPipelined[17]~67_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sReadCountPipelined_0),
	.q(\sReadCountPipelined[17]~q ),
	.prn(vcc));
defparam \sReadCountPipelined[17] .is_wysiwyg = "true";
defparam \sReadCountPipelined[17] .power_up = "low";

cycloneive_lcell_comb \sReadCountPipelined[18]~69 (
	.dataa(\sReadCountPipelined[18]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCountPipelined[17]~68 ),
	.combout(\sReadCountPipelined[18]~69_combout ),
	.cout(\sReadCountPipelined[18]~70 ));
defparam \sReadCountPipelined[18]~69 .lut_mask = 16'h5AAF;
defparam \sReadCountPipelined[18]~69 .sum_lutc_input = "cin";

dffeas \sReadCountPipelined[18] (
	.clk(Clk),
	.d(\sReadCountPipelined[18]~69_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sReadCountPipelined_0),
	.q(\sReadCountPipelined[18]~q ),
	.prn(vcc));
defparam \sReadCountPipelined[18] .is_wysiwyg = "true";
defparam \sReadCountPipelined[18] .power_up = "low";

cycloneive_lcell_comb \sReadCountPipelined[19]~71 (
	.dataa(\sReadCountPipelined[19]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCountPipelined[18]~70 ),
	.combout(\sReadCountPipelined[19]~71_combout ),
	.cout(\sReadCountPipelined[19]~72 ));
defparam \sReadCountPipelined[19]~71 .lut_mask = 16'h5A5F;
defparam \sReadCountPipelined[19]~71 .sum_lutc_input = "cin";

dffeas \sReadCountPipelined[19] (
	.clk(Clk),
	.d(\sReadCountPipelined[19]~71_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sReadCountPipelined_0),
	.q(\sReadCountPipelined[19]~q ),
	.prn(vcc));
defparam \sReadCountPipelined[19] .is_wysiwyg = "true";
defparam \sReadCountPipelined[19] .power_up = "low";

cycloneive_lcell_comb \sReadCountPipelined[20]~73 (
	.dataa(\sReadCountPipelined[20]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCountPipelined[19]~72 ),
	.combout(\sReadCountPipelined[20]~73_combout ),
	.cout(\sReadCountPipelined[20]~74 ));
defparam \sReadCountPipelined[20]~73 .lut_mask = 16'h5AAF;
defparam \sReadCountPipelined[20]~73 .sum_lutc_input = "cin";

dffeas \sReadCountPipelined[20] (
	.clk(Clk),
	.d(\sReadCountPipelined[20]~73_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sReadCountPipelined_0),
	.q(\sReadCountPipelined[20]~q ),
	.prn(vcc));
defparam \sReadCountPipelined[20] .is_wysiwyg = "true";
defparam \sReadCountPipelined[20] .power_up = "low";

dffeas \sRegByteEnable[19] (
	.clk(Clk),
	.d(d_writedata_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sRegByteEnable[16]~4_combout ),
	.q(\sRegByteEnable[19]~q ),
	.prn(vcc));
defparam \sRegByteEnable[19] .is_wysiwyg = "true";
defparam \sRegByteEnable[19] .power_up = "low";

dffeas \sReg[19] (
	.clk(Clk),
	.d(d_writedata_19),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReg[0]~0_combout ),
	.q(\sReg[19]~q ),
	.prn(vcc));
defparam \sReg[19] .is_wysiwyg = "true";
defparam \sReg[19] .power_up = "low";

cycloneive_lcell_comb \ReadData[19]~36 (
	.dataa(W_alu_result_3),
	.datab(\sRegByteEnable[19]~q ),
	.datac(W_alu_result_2),
	.datad(\sReg[19]~q ),
	.cin(gnd),
	.combout(\ReadData[19]~36_combout ),
	.cout());
defparam \ReadData[19]~36 .lut_mask = 16'hFFDE;
defparam \ReadData[19]~36 .sum_lutc_input = "datac";

dffeas \sRegByteEnable[18] (
	.clk(Clk),
	.d(d_writedata_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sRegByteEnable[16]~4_combout ),
	.q(\sRegByteEnable[18]~q ),
	.prn(vcc));
defparam \sRegByteEnable[18] .is_wysiwyg = "true";
defparam \sRegByteEnable[18] .power_up = "low";

dffeas \sReg[18] (
	.clk(Clk),
	.d(d_writedata_18),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReg[0]~0_combout ),
	.q(\sReg[18]~q ),
	.prn(vcc));
defparam \sReg[18] .is_wysiwyg = "true";
defparam \sReg[18] .power_up = "low";

cycloneive_lcell_comb \ReadData[18]~38 (
	.dataa(W_alu_result_2),
	.datab(\sReadCount[18]~q ),
	.datac(W_alu_result_3),
	.datad(\sReg[18]~q ),
	.cin(gnd),
	.combout(\ReadData[18]~38_combout ),
	.cout());
defparam \ReadData[18]~38 .lut_mask = 16'hFFDE;
defparam \ReadData[18]~38 .sum_lutc_input = "datac";

dffeas \sRegByteEnable[17] (
	.clk(Clk),
	.d(d_writedata_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sRegByteEnable[16]~4_combout ),
	.q(\sRegByteEnable[17]~q ),
	.prn(vcc));
defparam \sRegByteEnable[17] .is_wysiwyg = "true";
defparam \sRegByteEnable[17] .power_up = "low";

dffeas \sReg[17] (
	.clk(Clk),
	.d(d_writedata_17),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReg[0]~0_combout ),
	.q(\sReg[17]~q ),
	.prn(vcc));
defparam \sReg[17] .is_wysiwyg = "true";
defparam \sReg[17] .power_up = "low";

cycloneive_lcell_comb \ReadData[17]~40 (
	.dataa(W_alu_result_3),
	.datab(\sRegByteEnable[17]~q ),
	.datac(W_alu_result_2),
	.datad(\sReg[17]~q ),
	.cin(gnd),
	.combout(\ReadData[17]~40_combout ),
	.cout());
defparam \ReadData[17]~40 .lut_mask = 16'hFFDE;
defparam \ReadData[17]~40 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sReadCount[21]~75 (
	.dataa(\sReadCount[21]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCount[20]~74 ),
	.combout(\sReadCount[21]~75_combout ),
	.cout(\sReadCount[21]~76 ));
defparam \sReadCount[21]~75 .lut_mask = 16'h5A5F;
defparam \sReadCount[21]~75 .sum_lutc_input = "cin";

dffeas \sReadCount[21] (
	.clk(Clk),
	.d(\sReadCount[21]~75_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReadCount[0]~34_combout ),
	.q(\sReadCount[21]~q ),
	.prn(vcc));
defparam \sReadCount[21] .is_wysiwyg = "true";
defparam \sReadCount[21] .power_up = "low";

cycloneive_lcell_comb \sReadCount[22]~77 (
	.dataa(\sReadCount[22]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCount[21]~76 ),
	.combout(\sReadCount[22]~77_combout ),
	.cout(\sReadCount[22]~78 ));
defparam \sReadCount[22]~77 .lut_mask = 16'h5AAF;
defparam \sReadCount[22]~77 .sum_lutc_input = "cin";

dffeas \sReadCount[22] (
	.clk(Clk),
	.d(\sReadCount[22]~77_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReadCount[0]~34_combout ),
	.q(\sReadCount[22]~q ),
	.prn(vcc));
defparam \sReadCount[22] .is_wysiwyg = "true";
defparam \sReadCount[22] .power_up = "low";

cycloneive_lcell_comb \sReadCount[23]~79 (
	.dataa(\sReadCount[23]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCount[22]~78 ),
	.combout(\sReadCount[23]~79_combout ),
	.cout(\sReadCount[23]~80 ));
defparam \sReadCount[23]~79 .lut_mask = 16'h5A5F;
defparam \sReadCount[23]~79 .sum_lutc_input = "cin";

dffeas \sReadCount[23] (
	.clk(Clk),
	.d(\sReadCount[23]~79_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReadCount[0]~34_combout ),
	.q(\sReadCount[23]~q ),
	.prn(vcc));
defparam \sReadCount[23] .is_wysiwyg = "true";
defparam \sReadCount[23] .power_up = "low";

dffeas \sRegByteEnable[23] (
	.clk(Clk),
	.d(d_writedata_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sRegByteEnable[16]~4_combout ),
	.q(\sRegByteEnable[23]~q ),
	.prn(vcc));
defparam \sRegByteEnable[23] .is_wysiwyg = "true";
defparam \sRegByteEnable[23] .power_up = "low";

dffeas \sReg[23] (
	.clk(Clk),
	.d(d_writedata_23),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReg[0]~0_combout ),
	.q(\sReg[23]~q ),
	.prn(vcc));
defparam \sReg[23] .is_wysiwyg = "true";
defparam \sReg[23] .power_up = "low";

cycloneive_lcell_comb \ReadData[23]~42 (
	.dataa(W_alu_result_3),
	.datab(\sRegByteEnable[23]~q ),
	.datac(W_alu_result_2),
	.datad(\sReg[23]~q ),
	.cin(gnd),
	.combout(\ReadData[23]~42_combout ),
	.cout());
defparam \ReadData[23]~42 .lut_mask = 16'hFFDE;
defparam \ReadData[23]~42 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sReadCountPipelined[21]~75 (
	.dataa(\sReadCountPipelined[21]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCountPipelined[20]~74 ),
	.combout(\sReadCountPipelined[21]~75_combout ),
	.cout(\sReadCountPipelined[21]~76 ));
defparam \sReadCountPipelined[21]~75 .lut_mask = 16'h5A5F;
defparam \sReadCountPipelined[21]~75 .sum_lutc_input = "cin";

dffeas \sReadCountPipelined[21] (
	.clk(Clk),
	.d(\sReadCountPipelined[21]~75_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sReadCountPipelined_0),
	.q(\sReadCountPipelined[21]~q ),
	.prn(vcc));
defparam \sReadCountPipelined[21] .is_wysiwyg = "true";
defparam \sReadCountPipelined[21] .power_up = "low";

cycloneive_lcell_comb \sReadCountPipelined[22]~77 (
	.dataa(\sReadCountPipelined[22]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCountPipelined[21]~76 ),
	.combout(\sReadCountPipelined[22]~77_combout ),
	.cout(\sReadCountPipelined[22]~78 ));
defparam \sReadCountPipelined[22]~77 .lut_mask = 16'h5AAF;
defparam \sReadCountPipelined[22]~77 .sum_lutc_input = "cin";

dffeas \sReadCountPipelined[22] (
	.clk(Clk),
	.d(\sReadCountPipelined[22]~77_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sReadCountPipelined_0),
	.q(\sReadCountPipelined[22]~q ),
	.prn(vcc));
defparam \sReadCountPipelined[22] .is_wysiwyg = "true";
defparam \sReadCountPipelined[22] .power_up = "low";

cycloneive_lcell_comb \sReadCountPipelined[23]~79 (
	.dataa(\sReadCountPipelined[23]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCountPipelined[22]~78 ),
	.combout(\sReadCountPipelined[23]~79_combout ),
	.cout(\sReadCountPipelined[23]~80 ));
defparam \sReadCountPipelined[23]~79 .lut_mask = 16'h5A5F;
defparam \sReadCountPipelined[23]~79 .sum_lutc_input = "cin";

dffeas \sReadCountPipelined[23] (
	.clk(Clk),
	.d(\sReadCountPipelined[23]~79_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sReadCountPipelined_0),
	.q(\sReadCountPipelined[23]~q ),
	.prn(vcc));
defparam \sReadCountPipelined[23] .is_wysiwyg = "true";
defparam \sReadCountPipelined[23] .power_up = "low";

dffeas \sRegByteEnable[22] (
	.clk(Clk),
	.d(d_writedata_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sRegByteEnable[16]~4_combout ),
	.q(\sRegByteEnable[22]~q ),
	.prn(vcc));
defparam \sRegByteEnable[22] .is_wysiwyg = "true";
defparam \sRegByteEnable[22] .power_up = "low";

dffeas \sReg[22] (
	.clk(Clk),
	.d(d_writedata_22),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReg[0]~0_combout ),
	.q(\sReg[22]~q ),
	.prn(vcc));
defparam \sReg[22] .is_wysiwyg = "true";
defparam \sReg[22] .power_up = "low";

cycloneive_lcell_comb \ReadData[22]~44 (
	.dataa(W_alu_result_2),
	.datab(\sReadCount[22]~q ),
	.datac(W_alu_result_3),
	.datad(\sReg[22]~q ),
	.cin(gnd),
	.combout(\ReadData[22]~44_combout ),
	.cout());
defparam \ReadData[22]~44 .lut_mask = 16'hFFDE;
defparam \ReadData[22]~44 .sum_lutc_input = "datac";

dffeas \sRegByteEnable[21] (
	.clk(Clk),
	.d(d_writedata_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sRegByteEnable[16]~4_combout ),
	.q(\sRegByteEnable[21]~q ),
	.prn(vcc));
defparam \sRegByteEnable[21] .is_wysiwyg = "true";
defparam \sRegByteEnable[21] .power_up = "low";

dffeas \sReg[21] (
	.clk(Clk),
	.d(d_writedata_21),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReg[0]~0_combout ),
	.q(\sReg[21]~q ),
	.prn(vcc));
defparam \sReg[21] .is_wysiwyg = "true";
defparam \sReg[21] .power_up = "low";

cycloneive_lcell_comb \ReadData[21]~46 (
	.dataa(W_alu_result_3),
	.datab(\sRegByteEnable[21]~q ),
	.datac(W_alu_result_2),
	.datad(\sReg[21]~q ),
	.cin(gnd),
	.combout(\ReadData[21]~46_combout ),
	.cout());
defparam \ReadData[21]~46 .lut_mask = 16'hFFDE;
defparam \ReadData[21]~46 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sRegByteEnable[24]~5 (
	.dataa(d_byteenable_3),
	.datab(\sRegByteEnable[24]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sRegByteEnable[24]~5_combout ),
	.cout());
defparam \sRegByteEnable[24]~5 .lut_mask = 16'hEEEE;
defparam \sRegByteEnable[24]~5 .sum_lutc_input = "datac";

dffeas \sRegByteEnable[24] (
	.clk(Clk),
	.d(d_writedata_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sRegByteEnable[24]~5_combout ),
	.q(\sRegByteEnable[24]~q ),
	.prn(vcc));
defparam \sRegByteEnable[24] .is_wysiwyg = "true";
defparam \sRegByteEnable[24] .power_up = "low";

cycloneive_lcell_comb \sReadCount[24]~81 (
	.dataa(\sReadCount[24]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCount[23]~80 ),
	.combout(\sReadCount[24]~81_combout ),
	.cout(\sReadCount[24]~82 ));
defparam \sReadCount[24]~81 .lut_mask = 16'h5AAF;
defparam \sReadCount[24]~81 .sum_lutc_input = "cin";

dffeas \sReadCount[24] (
	.clk(Clk),
	.d(\sReadCount[24]~81_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReadCount[0]~34_combout ),
	.q(\sReadCount[24]~q ),
	.prn(vcc));
defparam \sReadCount[24] .is_wysiwyg = "true";
defparam \sReadCount[24] .power_up = "low";

dffeas \sReg[24] (
	.clk(Clk),
	.d(d_writedata_24),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReg[0]~0_combout ),
	.q(\sReg[24]~q ),
	.prn(vcc));
defparam \sReg[24] .is_wysiwyg = "true";
defparam \sReg[24] .power_up = "low";

cycloneive_lcell_comb \ReadData[24]~48 (
	.dataa(W_alu_result_2),
	.datab(\sReadCount[24]~q ),
	.datac(W_alu_result_3),
	.datad(\sReg[24]~q ),
	.cin(gnd),
	.combout(\ReadData[24]~48_combout ),
	.cout());
defparam \ReadData[24]~48 .lut_mask = 16'hFFDE;
defparam \ReadData[24]~48 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sReadCountPipelined[24]~81 (
	.dataa(\sReadCountPipelined[24]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCountPipelined[23]~80 ),
	.combout(\sReadCountPipelined[24]~81_combout ),
	.cout(\sReadCountPipelined[24]~82 ));
defparam \sReadCountPipelined[24]~81 .lut_mask = 16'h5AAF;
defparam \sReadCountPipelined[24]~81 .sum_lutc_input = "cin";

dffeas \sReadCountPipelined[24] (
	.clk(Clk),
	.d(\sReadCountPipelined[24]~81_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sReadCountPipelined_0),
	.q(\sReadCountPipelined[24]~q ),
	.prn(vcc));
defparam \sReadCountPipelined[24] .is_wysiwyg = "true";
defparam \sReadCountPipelined[24] .power_up = "low";

cycloneive_lcell_comb \sReadCount[25]~83 (
	.dataa(\sReadCount[25]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCount[24]~82 ),
	.combout(\sReadCount[25]~83_combout ),
	.cout(\sReadCount[25]~84 ));
defparam \sReadCount[25]~83 .lut_mask = 16'h5A5F;
defparam \sReadCount[25]~83 .sum_lutc_input = "cin";

dffeas \sReadCount[25] (
	.clk(Clk),
	.d(\sReadCount[25]~83_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReadCount[0]~34_combout ),
	.q(\sReadCount[25]~q ),
	.prn(vcc));
defparam \sReadCount[25] .is_wysiwyg = "true";
defparam \sReadCount[25] .power_up = "low";

cycloneive_lcell_comb \sReadCount[26]~85 (
	.dataa(\sReadCount[26]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCount[25]~84 ),
	.combout(\sReadCount[26]~85_combout ),
	.cout(\sReadCount[26]~86 ));
defparam \sReadCount[26]~85 .lut_mask = 16'h5AAF;
defparam \sReadCount[26]~85 .sum_lutc_input = "cin";

dffeas \sReadCount[26] (
	.clk(Clk),
	.d(\sReadCount[26]~85_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReadCount[0]~34_combout ),
	.q(\sReadCount[26]~q ),
	.prn(vcc));
defparam \sReadCount[26] .is_wysiwyg = "true";
defparam \sReadCount[26] .power_up = "low";

cycloneive_lcell_comb \sReadCount[27]~87 (
	.dataa(\sReadCount[27]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCount[26]~86 ),
	.combout(\sReadCount[27]~87_combout ),
	.cout(\sReadCount[27]~88 ));
defparam \sReadCount[27]~87 .lut_mask = 16'h5A5F;
defparam \sReadCount[27]~87 .sum_lutc_input = "cin";

dffeas \sReadCount[27] (
	.clk(Clk),
	.d(\sReadCount[27]~87_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReadCount[0]~34_combout ),
	.q(\sReadCount[27]~q ),
	.prn(vcc));
defparam \sReadCount[27] .is_wysiwyg = "true";
defparam \sReadCount[27] .power_up = "low";

cycloneive_lcell_comb \sReadCount[28]~89 (
	.dataa(\sReadCount[28]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCount[27]~88 ),
	.combout(\sReadCount[28]~89_combout ),
	.cout(\sReadCount[28]~90 ));
defparam \sReadCount[28]~89 .lut_mask = 16'h5AAF;
defparam \sReadCount[28]~89 .sum_lutc_input = "cin";

dffeas \sReadCount[28] (
	.clk(Clk),
	.d(\sReadCount[28]~89_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReadCount[0]~34_combout ),
	.q(\sReadCount[28]~q ),
	.prn(vcc));
defparam \sReadCount[28] .is_wysiwyg = "true";
defparam \sReadCount[28] .power_up = "low";

cycloneive_lcell_comb \sReadCount[29]~91 (
	.dataa(\sReadCount[29]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCount[28]~90 ),
	.combout(\sReadCount[29]~91_combout ),
	.cout(\sReadCount[29]~92 ));
defparam \sReadCount[29]~91 .lut_mask = 16'h5A5F;
defparam \sReadCount[29]~91 .sum_lutc_input = "cin";

dffeas \sReadCount[29] (
	.clk(Clk),
	.d(\sReadCount[29]~91_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReadCount[0]~34_combout ),
	.q(\sReadCount[29]~q ),
	.prn(vcc));
defparam \sReadCount[29] .is_wysiwyg = "true";
defparam \sReadCount[29] .power_up = "low";

cycloneive_lcell_comb \sReadCount[30]~93 (
	.dataa(\sReadCount[30]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCount[29]~92 ),
	.combout(\sReadCount[30]~93_combout ),
	.cout(\sReadCount[30]~94 ));
defparam \sReadCount[30]~93 .lut_mask = 16'h5AAF;
defparam \sReadCount[30]~93 .sum_lutc_input = "cin";

dffeas \sReadCount[30] (
	.clk(Clk),
	.d(\sReadCount[30]~93_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReadCount[0]~34_combout ),
	.q(\sReadCount[30]~q ),
	.prn(vcc));
defparam \sReadCount[30] .is_wysiwyg = "true";
defparam \sReadCount[30] .power_up = "low";

cycloneive_lcell_comb \sReadCount[31]~95 (
	.dataa(\sReadCount[31]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\sReadCount[30]~94 ),
	.combout(\sReadCount[31]~95_combout ),
	.cout());
defparam \sReadCount[31]~95 .lut_mask = 16'h5A5A;
defparam \sReadCount[31]~95 .sum_lutc_input = "cin";

dffeas \sReadCount[31] (
	.clk(Clk),
	.d(\sReadCount[31]~95_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReadCount[0]~34_combout ),
	.q(\sReadCount[31]~q ),
	.prn(vcc));
defparam \sReadCount[31] .is_wysiwyg = "true";
defparam \sReadCount[31] .power_up = "low";

dffeas \sRegByteEnable[31] (
	.clk(Clk),
	.d(d_writedata_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sRegByteEnable[24]~5_combout ),
	.q(\sRegByteEnable[31]~q ),
	.prn(vcc));
defparam \sRegByteEnable[31] .is_wysiwyg = "true";
defparam \sRegByteEnable[31] .power_up = "low";

dffeas \sReg[31] (
	.clk(Clk),
	.d(d_writedata_31),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReg[0]~0_combout ),
	.q(\sReg[31]~q ),
	.prn(vcc));
defparam \sReg[31] .is_wysiwyg = "true";
defparam \sReg[31] .power_up = "low";

cycloneive_lcell_comb \ReadData[31]~50 (
	.dataa(W_alu_result_3),
	.datab(\sRegByteEnable[31]~q ),
	.datac(W_alu_result_2),
	.datad(\sReg[31]~q ),
	.cin(gnd),
	.combout(\ReadData[31]~50_combout ),
	.cout());
defparam \ReadData[31]~50 .lut_mask = 16'hFFDE;
defparam \ReadData[31]~50 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sReadCountPipelined[25]~83 (
	.dataa(\sReadCountPipelined[25]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCountPipelined[24]~82 ),
	.combout(\sReadCountPipelined[25]~83_combout ),
	.cout(\sReadCountPipelined[25]~84 ));
defparam \sReadCountPipelined[25]~83 .lut_mask = 16'h5A5F;
defparam \sReadCountPipelined[25]~83 .sum_lutc_input = "cin";

dffeas \sReadCountPipelined[25] (
	.clk(Clk),
	.d(\sReadCountPipelined[25]~83_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sReadCountPipelined_0),
	.q(\sReadCountPipelined[25]~q ),
	.prn(vcc));
defparam \sReadCountPipelined[25] .is_wysiwyg = "true";
defparam \sReadCountPipelined[25] .power_up = "low";

cycloneive_lcell_comb \sReadCountPipelined[26]~85 (
	.dataa(\sReadCountPipelined[26]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCountPipelined[25]~84 ),
	.combout(\sReadCountPipelined[26]~85_combout ),
	.cout(\sReadCountPipelined[26]~86 ));
defparam \sReadCountPipelined[26]~85 .lut_mask = 16'h5AAF;
defparam \sReadCountPipelined[26]~85 .sum_lutc_input = "cin";

dffeas \sReadCountPipelined[26] (
	.clk(Clk),
	.d(\sReadCountPipelined[26]~85_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sReadCountPipelined_0),
	.q(\sReadCountPipelined[26]~q ),
	.prn(vcc));
defparam \sReadCountPipelined[26] .is_wysiwyg = "true";
defparam \sReadCountPipelined[26] .power_up = "low";

cycloneive_lcell_comb \sReadCountPipelined[27]~87 (
	.dataa(\sReadCountPipelined[27]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCountPipelined[26]~86 ),
	.combout(\sReadCountPipelined[27]~87_combout ),
	.cout(\sReadCountPipelined[27]~88 ));
defparam \sReadCountPipelined[27]~87 .lut_mask = 16'h5A5F;
defparam \sReadCountPipelined[27]~87 .sum_lutc_input = "cin";

dffeas \sReadCountPipelined[27] (
	.clk(Clk),
	.d(\sReadCountPipelined[27]~87_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sReadCountPipelined_0),
	.q(\sReadCountPipelined[27]~q ),
	.prn(vcc));
defparam \sReadCountPipelined[27] .is_wysiwyg = "true";
defparam \sReadCountPipelined[27] .power_up = "low";

cycloneive_lcell_comb \sReadCountPipelined[28]~89 (
	.dataa(\sReadCountPipelined[28]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCountPipelined[27]~88 ),
	.combout(\sReadCountPipelined[28]~89_combout ),
	.cout(\sReadCountPipelined[28]~90 ));
defparam \sReadCountPipelined[28]~89 .lut_mask = 16'h5AAF;
defparam \sReadCountPipelined[28]~89 .sum_lutc_input = "cin";

dffeas \sReadCountPipelined[28] (
	.clk(Clk),
	.d(\sReadCountPipelined[28]~89_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sReadCountPipelined_0),
	.q(\sReadCountPipelined[28]~q ),
	.prn(vcc));
defparam \sReadCountPipelined[28] .is_wysiwyg = "true";
defparam \sReadCountPipelined[28] .power_up = "low";

cycloneive_lcell_comb \sReadCountPipelined[29]~91 (
	.dataa(\sReadCountPipelined[29]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCountPipelined[28]~90 ),
	.combout(\sReadCountPipelined[29]~91_combout ),
	.cout(\sReadCountPipelined[29]~92 ));
defparam \sReadCountPipelined[29]~91 .lut_mask = 16'h5A5F;
defparam \sReadCountPipelined[29]~91 .sum_lutc_input = "cin";

dffeas \sReadCountPipelined[29] (
	.clk(Clk),
	.d(\sReadCountPipelined[29]~91_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sReadCountPipelined_0),
	.q(\sReadCountPipelined[29]~q ),
	.prn(vcc));
defparam \sReadCountPipelined[29] .is_wysiwyg = "true";
defparam \sReadCountPipelined[29] .power_up = "low";

cycloneive_lcell_comb \sReadCountPipelined[30]~93 (
	.dataa(\sReadCountPipelined[30]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\sReadCountPipelined[29]~92 ),
	.combout(\sReadCountPipelined[30]~93_combout ),
	.cout(\sReadCountPipelined[30]~94 ));
defparam \sReadCountPipelined[30]~93 .lut_mask = 16'h5AAF;
defparam \sReadCountPipelined[30]~93 .sum_lutc_input = "cin";

dffeas \sReadCountPipelined[30] (
	.clk(Clk),
	.d(\sReadCountPipelined[30]~93_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sReadCountPipelined_0),
	.q(\sReadCountPipelined[30]~q ),
	.prn(vcc));
defparam \sReadCountPipelined[30] .is_wysiwyg = "true";
defparam \sReadCountPipelined[30] .power_up = "low";

cycloneive_lcell_comb \sReadCountPipelined[31]~95 (
	.dataa(\sReadCountPipelined[31]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\sReadCountPipelined[30]~94 ),
	.combout(\sReadCountPipelined[31]~95_combout ),
	.cout());
defparam \sReadCountPipelined[31]~95 .lut_mask = 16'h5A5A;
defparam \sReadCountPipelined[31]~95 .sum_lutc_input = "cin";

dffeas \sReadCountPipelined[31] (
	.clk(Clk),
	.d(\sReadCountPipelined[31]~95_combout ),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sReadCountPipelined_0),
	.q(\sReadCountPipelined[31]~q ),
	.prn(vcc));
defparam \sReadCountPipelined[31] .is_wysiwyg = "true";
defparam \sReadCountPipelined[31] .power_up = "low";

dffeas \sRegByteEnable[30] (
	.clk(Clk),
	.d(d_writedata_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sRegByteEnable[24]~5_combout ),
	.q(\sRegByteEnable[30]~q ),
	.prn(vcc));
defparam \sRegByteEnable[30] .is_wysiwyg = "true";
defparam \sRegByteEnable[30] .power_up = "low";

dffeas \sReg[30] (
	.clk(Clk),
	.d(d_writedata_30),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReg[0]~0_combout ),
	.q(\sReg[30]~q ),
	.prn(vcc));
defparam \sReg[30] .is_wysiwyg = "true";
defparam \sReg[30] .power_up = "low";

cycloneive_lcell_comb \ReadData[30]~52 (
	.dataa(W_alu_result_2),
	.datab(\sReadCount[30]~q ),
	.datac(W_alu_result_3),
	.datad(\sReg[30]~q ),
	.cin(gnd),
	.combout(\ReadData[30]~52_combout ),
	.cout());
defparam \ReadData[30]~52 .lut_mask = 16'hFFDE;
defparam \ReadData[30]~52 .sum_lutc_input = "datac";

dffeas \sRegByteEnable[29] (
	.clk(Clk),
	.d(d_writedata_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sRegByteEnable[24]~5_combout ),
	.q(\sRegByteEnable[29]~q ),
	.prn(vcc));
defparam \sRegByteEnable[29] .is_wysiwyg = "true";
defparam \sRegByteEnable[29] .power_up = "low";

dffeas \sReg[29] (
	.clk(Clk),
	.d(d_writedata_29),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReg[0]~0_combout ),
	.q(\sReg[29]~q ),
	.prn(vcc));
defparam \sReg[29] .is_wysiwyg = "true";
defparam \sReg[29] .power_up = "low";

cycloneive_lcell_comb \ReadData[29]~54 (
	.dataa(W_alu_result_3),
	.datab(\sRegByteEnable[29]~q ),
	.datac(W_alu_result_2),
	.datad(\sReg[29]~q ),
	.cin(gnd),
	.combout(\ReadData[29]~54_combout ),
	.cout());
defparam \ReadData[29]~54 .lut_mask = 16'hFFDE;
defparam \ReadData[29]~54 .sum_lutc_input = "datac";

dffeas \sRegByteEnable[28] (
	.clk(Clk),
	.d(d_writedata_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sRegByteEnable[24]~5_combout ),
	.q(\sRegByteEnable[28]~q ),
	.prn(vcc));
defparam \sRegByteEnable[28] .is_wysiwyg = "true";
defparam \sRegByteEnable[28] .power_up = "low";

dffeas \sReg[28] (
	.clk(Clk),
	.d(d_writedata_28),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReg[0]~0_combout ),
	.q(\sReg[28]~q ),
	.prn(vcc));
defparam \sReg[28] .is_wysiwyg = "true";
defparam \sReg[28] .power_up = "low";

cycloneive_lcell_comb \ReadData[28]~56 (
	.dataa(W_alu_result_2),
	.datab(\sReadCount[28]~q ),
	.datac(W_alu_result_3),
	.datad(\sReg[28]~q ),
	.cin(gnd),
	.combout(\ReadData[28]~56_combout ),
	.cout());
defparam \ReadData[28]~56 .lut_mask = 16'hFFDE;
defparam \ReadData[28]~56 .sum_lutc_input = "datac";

dffeas \sRegByteEnable[27] (
	.clk(Clk),
	.d(d_writedata_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sRegByteEnable[24]~5_combout ),
	.q(\sRegByteEnable[27]~q ),
	.prn(vcc));
defparam \sRegByteEnable[27] .is_wysiwyg = "true";
defparam \sRegByteEnable[27] .power_up = "low";

dffeas \sReg[27] (
	.clk(Clk),
	.d(d_writedata_27),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReg[0]~0_combout ),
	.q(\sReg[27]~q ),
	.prn(vcc));
defparam \sReg[27] .is_wysiwyg = "true";
defparam \sReg[27] .power_up = "low";

cycloneive_lcell_comb \ReadData[27]~58 (
	.dataa(W_alu_result_3),
	.datab(\sRegByteEnable[27]~q ),
	.datac(W_alu_result_2),
	.datad(\sReg[27]~q ),
	.cin(gnd),
	.combout(\ReadData[27]~58_combout ),
	.cout());
defparam \ReadData[27]~58 .lut_mask = 16'hFFDE;
defparam \ReadData[27]~58 .sum_lutc_input = "datac";

dffeas \sRegByteEnable[26] (
	.clk(Clk),
	.d(d_writedata_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sRegByteEnable[24]~5_combout ),
	.q(\sRegByteEnable[26]~q ),
	.prn(vcc));
defparam \sRegByteEnable[26] .is_wysiwyg = "true";
defparam \sRegByteEnable[26] .power_up = "low";

dffeas \sReg[26] (
	.clk(Clk),
	.d(d_writedata_26),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReg[0]~0_combout ),
	.q(\sReg[26]~q ),
	.prn(vcc));
defparam \sReg[26] .is_wysiwyg = "true";
defparam \sReg[26] .power_up = "low";

cycloneive_lcell_comb \ReadData[26]~60 (
	.dataa(W_alu_result_2),
	.datab(\sReadCount[26]~q ),
	.datac(W_alu_result_3),
	.datad(\sReg[26]~q ),
	.cin(gnd),
	.combout(\ReadData[26]~60_combout ),
	.cout());
defparam \ReadData[26]~60 .lut_mask = 16'hFFDE;
defparam \ReadData[26]~60 .sum_lutc_input = "datac";

dffeas \sRegByteEnable[25] (
	.clk(Clk),
	.d(d_writedata_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sRegByteEnable[24]~5_combout ),
	.q(\sRegByteEnable[25]~q ),
	.prn(vcc));
defparam \sRegByteEnable[25] .is_wysiwyg = "true";
defparam \sRegByteEnable[25] .power_up = "low";

dffeas \sReg[25] (
	.clk(Clk),
	.d(d_writedata_25),
	.asdata(vcc),
	.clrn(Reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sReg[0]~0_combout ),
	.q(\sReg[25]~q ),
	.prn(vcc));
defparam \sReg[25] .is_wysiwyg = "true";
defparam \sReg[25] .power_up = "low";

cycloneive_lcell_comb \ReadData[25]~62 (
	.dataa(W_alu_result_3),
	.datab(\sRegByteEnable[25]~q ),
	.datac(W_alu_result_2),
	.datad(\sReg[25]~q ),
	.cin(gnd),
	.combout(\ReadData[25]~62_combout ),
	.cout());
defparam \ReadData[25]~62 .lut_mask = 16'hFFDE;
defparam \ReadData[25]~62 .sum_lutc_input = "datac";

endmodule

module nios_mcu_nios_mcu_jtag_uart_0 (
	W_alu_result_2,
	adapted_tdo,
	d_writedata_0,
	r_sync_rst,
	rst1,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	read_latency_shift_reg,
	m0_write,
	Equal3,
	av_waitrequest1,
	mem_used_1,
	always2,
	b_full,
	read_01,
	av_readdata_0,
	av_readdata_9,
	av_readdata_8,
	d_writedata_10,
	av_readdata_1,
	av_readdata_2,
	av_readdata_3,
	av_readdata_4,
	av_readdata_5,
	av_readdata_6,
	av_readdata_7,
	b_non_empty,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_31,
	counter_reg_bit_01,
	counter_reg_bit_21,
	counter_reg_bit_11,
	b_full1,
	counter_reg_bit_51,
	counter_reg_bit_41,
	ac1,
	rvalid1,
	woverflow1,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	splitter_nodes_receive_0_3,
	virtual_ir_scan_reg,
	clr_reg,
	state_3,
	state_8,
	irf_reg_0_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_2;
output 	adapted_tdo;
input 	d_writedata_0;
input 	r_sync_rst;
output 	rst1;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	d_writedata_6;
input 	d_writedata_7;
input 	read_latency_shift_reg;
input 	m0_write;
input 	Equal3;
output 	av_waitrequest1;
input 	mem_used_1;
input 	always2;
output 	b_full;
output 	read_01;
output 	av_readdata_0;
output 	av_readdata_9;
output 	av_readdata_8;
input 	d_writedata_10;
output 	av_readdata_1;
output 	av_readdata_2;
output 	av_readdata_3;
output 	av_readdata_4;
output 	av_readdata_5;
output 	av_readdata_6;
output 	av_readdata_7;
output 	b_non_empty;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_31;
output 	counter_reg_bit_01;
output 	counter_reg_bit_21;
output 	counter_reg_bit_11;
output 	b_full1;
output 	counter_reg_bit_51;
output 	counter_reg_bit_41;
output 	ac1;
output 	rvalid1;
output 	woverflow1;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	splitter_nodes_receive_0_3;
input 	virtual_ir_scan_reg;
input 	clr_reg;
input 	state_3;
input 	state_8;
input 	irf_reg_0_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \t_dav~q ;
wire \nios_mcu_jtag_uart_0_alt_jtag_atlantic|rvalid0~q ;
wire \r_val~q ;
wire \nios_mcu_jtag_uart_0_alt_jtag_atlantic|r_ena1~q ;
wire \nios_mcu_jtag_uart_0_alt_jtag_atlantic|t_ena~reg0_q ;
wire \fifo_rd~0_combout ;
wire \the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ;
wire \r_val~0_combout ;
wire \fifo_wr~q ;
wire \wr_rfifo~combout ;
wire \nios_mcu_jtag_uart_0_alt_jtag_atlantic|wdata[0]~q ;
wire \nios_mcu_jtag_uart_0_alt_jtag_atlantic|t_pause~reg0_q ;
wire \nios_mcu_jtag_uart_0_alt_jtag_atlantic|wdata[1]~q ;
wire \nios_mcu_jtag_uart_0_alt_jtag_atlantic|wdata[2]~q ;
wire \nios_mcu_jtag_uart_0_alt_jtag_atlantic|wdata[3]~q ;
wire \nios_mcu_jtag_uart_0_alt_jtag_atlantic|wdata[4]~q ;
wire \nios_mcu_jtag_uart_0_alt_jtag_atlantic|wdata[5]~q ;
wire \nios_mcu_jtag_uart_0_alt_jtag_atlantic|wdata[6]~q ;
wire \nios_mcu_jtag_uart_0_alt_jtag_atlantic|wdata[7]~q ;
wire \fifo_wr~0_combout ;
wire \av_waitrequest~0_combout ;
wire \av_waitrequest~1_combout ;
wire \fifo_rd~1_combout ;
wire \ien_AE~0_combout ;
wire \ien_AF~q ;
wire \LessThan0~0_combout ;
wire \LessThan0~1_combout ;
wire \fifo_AE~q ;
wire \ien_AE~q ;
wire \pause_irq~0_combout ;
wire \pause_irq~q ;
wire \Add0~1 ;
wire \Add0~3 ;
wire \Add0~4_combout ;
wire \Add0~0_combout ;
wire \Add0~2_combout ;
wire \LessThan1~0_combout ;
wire \Add0~5 ;
wire \Add0~6_combout ;
wire \Add0~7 ;
wire \Add0~8_combout ;
wire \LessThan1~1_combout ;
wire \Add0~9 ;
wire \Add0~10_combout ;
wire \Add0~11 ;
wire \Add0~12_combout ;
wire \LessThan1~2_combout ;
wire \fifo_AF~q ;
wire \ac~0_combout ;
wire \ac~1_combout ;
wire \rvalid~0_combout ;
wire \woverflow~0_combout ;
wire \woverflow~1_combout ;


nios_mcu_alt_jtag_atlantic nios_mcu_jtag_uart_0_alt_jtag_atlantic(
	.r_dat({\the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[7] ,\the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[6] ,\the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[5] ,
\the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[4] ,\the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[3] ,\the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[2] ,
\the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[1] ,\the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[0] }),
	.adapted_tdo1(adapted_tdo),
	.rst_n(r_sync_rst),
	.rst11(rst1),
	.t_dav(\t_dav~q ),
	.rvalid01(\nios_mcu_jtag_uart_0_alt_jtag_atlantic|rvalid0~q ),
	.r_val(\r_val~q ),
	.r_ena11(\nios_mcu_jtag_uart_0_alt_jtag_atlantic|r_ena1~q ),
	.t_ena(\nios_mcu_jtag_uart_0_alt_jtag_atlantic|t_ena~reg0_q ),
	.wdata_0(\nios_mcu_jtag_uart_0_alt_jtag_atlantic|wdata[0]~q ),
	.t_pause(\nios_mcu_jtag_uart_0_alt_jtag_atlantic|t_pause~reg0_q ),
	.wdata_1(\nios_mcu_jtag_uart_0_alt_jtag_atlantic|wdata[1]~q ),
	.wdata_2(\nios_mcu_jtag_uart_0_alt_jtag_atlantic|wdata[2]~q ),
	.wdata_3(\nios_mcu_jtag_uart_0_alt_jtag_atlantic|wdata[3]~q ),
	.wdata_4(\nios_mcu_jtag_uart_0_alt_jtag_atlantic|wdata[4]~q ),
	.wdata_5(\nios_mcu_jtag_uart_0_alt_jtag_atlantic|wdata[5]~q ),
	.wdata_6(\nios_mcu_jtag_uart_0_alt_jtag_atlantic|wdata[6]~q ),
	.wdata_7(\nios_mcu_jtag_uart_0_alt_jtag_atlantic|wdata[7]~q ),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_4(state_4),
	.splitter_nodes_receive_0_3(splitter_nodes_receive_0_3),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.clr_reg(clr_reg),
	.state_3(state_3),
	.state_8(state_8),
	.irf_reg_0_1(irf_reg_0_1),
	.clk(clk_clk));

nios_mcu_nios_mcu_jtag_uart_0_scfifo_r the_nios_mcu_jtag_uart_0_scfifo_r(
	.q_b_0(\the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.q_b_1(\the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.q_b_2(\the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.q_b_3(\the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.q_b_4(\the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.q_b_5(\the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.q_b_6(\the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.q_b_7(\the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.r_sync_rst(r_sync_rst),
	.b_full(b_full),
	.b_non_empty(b_non_empty),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.t_ena(\nios_mcu_jtag_uart_0_alt_jtag_atlantic|t_ena~reg0_q ),
	.fifo_rd(\fifo_rd~0_combout ),
	.wr_rfifo(\wr_rfifo~combout ),
	.wdata_0(\nios_mcu_jtag_uart_0_alt_jtag_atlantic|wdata[0]~q ),
	.fifo_rd1(\fifo_rd~1_combout ),
	.wdata_1(\nios_mcu_jtag_uart_0_alt_jtag_atlantic|wdata[1]~q ),
	.wdata_2(\nios_mcu_jtag_uart_0_alt_jtag_atlantic|wdata[2]~q ),
	.wdata_3(\nios_mcu_jtag_uart_0_alt_jtag_atlantic|wdata[3]~q ),
	.wdata_4(\nios_mcu_jtag_uart_0_alt_jtag_atlantic|wdata[4]~q ),
	.wdata_5(\nios_mcu_jtag_uart_0_alt_jtag_atlantic|wdata[5]~q ),
	.wdata_6(\nios_mcu_jtag_uart_0_alt_jtag_atlantic|wdata[6]~q ),
	.wdata_7(\nios_mcu_jtag_uart_0_alt_jtag_atlantic|wdata[7]~q ),
	.clk_clk(clk_clk));

nios_mcu_nios_mcu_jtag_uart_0_scfifo_w the_nios_mcu_jtag_uart_0_scfifo_w(
	.q_b_7(\the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.q_b_0(\the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.q_b_1(\the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.q_b_2(\the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.q_b_3(\the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.q_b_4(\the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.q_b_5(\the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.q_b_6(\the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.d_writedata_0(d_writedata_0),
	.r_sync_rst(r_sync_rst),
	.d_writedata_1(d_writedata_1),
	.d_writedata_2(d_writedata_2),
	.d_writedata_3(d_writedata_3),
	.d_writedata_4(d_writedata_4),
	.d_writedata_5(d_writedata_5),
	.d_writedata_6(d_writedata_6),
	.d_writedata_7(d_writedata_7),
	.b_non_empty(\the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.r_val(\r_val~0_combout ),
	.fifo_wr(\fifo_wr~q ),
	.counter_reg_bit_3(counter_reg_bit_31),
	.counter_reg_bit_0(counter_reg_bit_01),
	.counter_reg_bit_2(counter_reg_bit_21),
	.counter_reg_bit_1(counter_reg_bit_11),
	.b_full(b_full1),
	.counter_reg_bit_5(counter_reg_bit_51),
	.counter_reg_bit_4(counter_reg_bit_41),
	.clk_clk(clk_clk));

dffeas t_dav(
	.clk(clk_clk),
	.d(b_full),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\t_dav~q ),
	.prn(vcc));
defparam t_dav.is_wysiwyg = "true";
defparam t_dav.power_up = "low";

dffeas r_val(
	.clk(clk_clk),
	.d(\r_val~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_val~q ),
	.prn(vcc));
defparam r_val.is_wysiwyg = "true";
defparam r_val.power_up = "low";

cycloneive_lcell_comb \fifo_rd~0 (
	.dataa(read_latency_shift_reg),
	.datab(\av_waitrequest~0_combout ),
	.datac(b_non_empty),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\fifo_rd~0_combout ),
	.cout());
defparam \fifo_rd~0 .lut_mask = 16'hFEFF;
defparam \fifo_rd~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \r_val~0 (
	.dataa(\the_nios_mcu_jtag_uart_0_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.datab(\r_val~q ),
	.datac(\nios_mcu_jtag_uart_0_alt_jtag_atlantic|r_ena1~q ),
	.datad(\nios_mcu_jtag_uart_0_alt_jtag_atlantic|rvalid0~q ),
	.cin(gnd),
	.combout(\r_val~0_combout ),
	.cout());
defparam \r_val~0 .lut_mask = 16'hBFFF;
defparam \r_val~0 .sum_lutc_input = "datac";

dffeas fifo_wr(
	.clk(clk_clk),
	.d(\fifo_wr~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_wr~q ),
	.prn(vcc));
defparam fifo_wr.is_wysiwyg = "true";
defparam fifo_wr.power_up = "low";

cycloneive_lcell_comb wr_rfifo(
	.dataa(\nios_mcu_jtag_uart_0_alt_jtag_atlantic|t_ena~reg0_q ),
	.datab(gnd),
	.datac(gnd),
	.datad(b_full),
	.cin(gnd),
	.combout(\wr_rfifo~combout ),
	.cout());
defparam wr_rfifo.lut_mask = 16'hAAFF;
defparam wr_rfifo.sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_wr~0 (
	.dataa(b_full1),
	.datab(gnd),
	.datac(gnd),
	.datad(\woverflow~0_combout ),
	.cin(gnd),
	.combout(\fifo_wr~0_combout ),
	.cout());
defparam \fifo_wr~0 .lut_mask = 16'hFF55;
defparam \fifo_wr~0 .sum_lutc_input = "datac";

dffeas av_waitrequest(
	.clk(clk_clk),
	.d(\av_waitrequest~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_waitrequest1),
	.prn(vcc));
defparam av_waitrequest.is_wysiwyg = "true";
defparam av_waitrequest.power_up = "low";

dffeas read_0(
	.clk(clk_clk),
	.d(\fifo_rd~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_01),
	.prn(vcc));
defparam read_0.is_wysiwyg = "true";
defparam read_0.power_up = "low";

cycloneive_lcell_comb \av_readdata[0]~0 (
	.dataa(\the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.datab(\ien_AF~q ),
	.datac(gnd),
	.datad(read_01),
	.cin(gnd),
	.combout(av_readdata_0),
	.cout());
defparam \av_readdata[0]~0 .lut_mask = 16'hAACC;
defparam \av_readdata[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata[9] (
	.dataa(\fifo_AE~q ),
	.datab(\ien_AE~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_9),
	.cout());
defparam \av_readdata[9] .lut_mask = 16'hEEEE;
defparam \av_readdata[9] .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata[8]~1 (
	.dataa(\ien_AF~q ),
	.datab(\pause_irq~q ),
	.datac(\fifo_AF~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_8),
	.cout());
defparam \av_readdata[8]~1 .lut_mask = 16'hFEFE;
defparam \av_readdata[8]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata[1]~2 (
	.dataa(\the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.datab(\ien_AE~q ),
	.datac(gnd),
	.datad(read_01),
	.cin(gnd),
	.combout(av_readdata_1),
	.cout());
defparam \av_readdata[1]~2 .lut_mask = 16'hAACC;
defparam \av_readdata[1]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata[2]~3 (
	.dataa(read_01),
	.datab(\the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_2),
	.cout());
defparam \av_readdata[2]~3 .lut_mask = 16'hEEEE;
defparam \av_readdata[2]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata[3]~4 (
	.dataa(read_01),
	.datab(\the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_3),
	.cout());
defparam \av_readdata[3]~4 .lut_mask = 16'hEEEE;
defparam \av_readdata[3]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata[4]~5 (
	.dataa(read_01),
	.datab(\the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_4),
	.cout());
defparam \av_readdata[4]~5 .lut_mask = 16'hEEEE;
defparam \av_readdata[4]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata[5]~6 (
	.dataa(read_01),
	.datab(\the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_5),
	.cout());
defparam \av_readdata[5]~6 .lut_mask = 16'hEEEE;
defparam \av_readdata[5]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata[6]~7 (
	.dataa(read_01),
	.datab(\the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_6),
	.cout());
defparam \av_readdata[6]~7 .lut_mask = 16'hEEEE;
defparam \av_readdata[6]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata[7]~8 (
	.dataa(read_01),
	.datab(\the_nios_mcu_jtag_uart_0_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(av_readdata_7),
	.cout());
defparam \av_readdata[7]~8 .lut_mask = 16'hEEEE;
defparam \av_readdata[7]~8 .sum_lutc_input = "datac";

dffeas ac(
	.clk(clk_clk),
	.d(\ac~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ac1),
	.prn(vcc));
defparam ac.is_wysiwyg = "true";
defparam ac.power_up = "low";

dffeas rvalid(
	.clk(clk_clk),
	.d(\rvalid~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rvalid1),
	.prn(vcc));
defparam rvalid.is_wysiwyg = "true";
defparam rvalid.power_up = "low";

dffeas woverflow(
	.clk(clk_clk),
	.d(\woverflow~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(woverflow1),
	.prn(vcc));
defparam woverflow.is_wysiwyg = "true";
defparam woverflow.power_up = "low";

cycloneive_lcell_comb \av_waitrequest~0 (
	.dataa(Equal3),
	.datab(gnd),
	.datac(av_waitrequest1),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\av_waitrequest~0_combout ),
	.cout());
defparam \av_waitrequest~0 .lut_mask = 16'hAFFF;
defparam \av_waitrequest~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_waitrequest~1 (
	.dataa(rst1),
	.datab(always2),
	.datac(\av_waitrequest~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\av_waitrequest~1_combout ),
	.cout());
defparam \av_waitrequest~1 .lut_mask = 16'hFEFE;
defparam \av_waitrequest~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_rd~1 (
	.dataa(read_latency_shift_reg),
	.datab(\av_waitrequest~0_combout ),
	.datac(gnd),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\fifo_rd~1_combout ),
	.cout());
defparam \fifo_rd~1 .lut_mask = 16'hEEFF;
defparam \fifo_rd~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ien_AE~0 (
	.dataa(rst1),
	.datab(W_alu_result_2),
	.datac(m0_write),
	.datad(\av_waitrequest~0_combout ),
	.cin(gnd),
	.combout(\ien_AE~0_combout ),
	.cout());
defparam \ien_AE~0 .lut_mask = 16'hFFFE;
defparam \ien_AE~0 .sum_lutc_input = "datac";

dffeas ien_AF(
	.clk(clk_clk),
	.d(d_writedata_0),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ien_AE~0_combout ),
	.q(\ien_AF~q ),
	.prn(vcc));
defparam ien_AF.is_wysiwyg = "true";
defparam ien_AF.power_up = "low";

cycloneive_lcell_comb \LessThan0~0 (
	.dataa(counter_reg_bit_31),
	.datab(counter_reg_bit_01),
	.datac(counter_reg_bit_21),
	.datad(counter_reg_bit_11),
	.cin(gnd),
	.combout(\LessThan0~0_combout ),
	.cout());
defparam \LessThan0~0 .lut_mask = 16'hFFFE;
defparam \LessThan0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \LessThan0~1 (
	.dataa(\LessThan0~0_combout ),
	.datab(b_full1),
	.datac(counter_reg_bit_51),
	.datad(counter_reg_bit_41),
	.cin(gnd),
	.combout(\LessThan0~1_combout ),
	.cout());
defparam \LessThan0~1 .lut_mask = 16'h7FFF;
defparam \LessThan0~1 .sum_lutc_input = "datac";

dffeas fifo_AE(
	.clk(clk_clk),
	.d(\LessThan0~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_AE~q ),
	.prn(vcc));
defparam fifo_AE.is_wysiwyg = "true";
defparam fifo_AE.power_up = "low";

dffeas ien_AE(
	.clk(clk_clk),
	.d(d_writedata_1),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ien_AE~0_combout ),
	.q(\ien_AE~q ),
	.prn(vcc));
defparam ien_AE.is_wysiwyg = "true";
defparam ien_AE.power_up = "low";

cycloneive_lcell_comb \pause_irq~0 (
	.dataa(b_non_empty),
	.datab(\nios_mcu_jtag_uart_0_alt_jtag_atlantic|t_pause~reg0_q ),
	.datac(\pause_irq~q ),
	.datad(read_01),
	.cin(gnd),
	.combout(\pause_irq~0_combout ),
	.cout());
defparam \pause_irq~0 .lut_mask = 16'hFEFF;
defparam \pause_irq~0 .sum_lutc_input = "datac";

dffeas pause_irq(
	.clk(clk_clk),
	.d(\pause_irq~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pause_irq~q ),
	.prn(vcc));
defparam pause_irq.is_wysiwyg = "true";
defparam pause_irq.power_up = "low";

cycloneive_lcell_comb \Add0~0 (
	.dataa(counter_reg_bit_0),
	.datab(counter_reg_bit_1),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout(\Add0~1 ));
defparam \Add0~0 .lut_mask = 16'h6677;
defparam \Add0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add0~2 (
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~1 ),
	.combout(\Add0~2_combout ),
	.cout(\Add0~3 ));
defparam \Add0~2 .lut_mask = 16'h5AAF;
defparam \Add0~2 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add0~4 (
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~3 ),
	.combout(\Add0~4_combout ),
	.cout(\Add0~5 ));
defparam \Add0~4 .lut_mask = 16'h5A5F;
defparam \Add0~4 .sum_lutc_input = "cin";

cycloneive_lcell_comb \LessThan1~0 (
	.dataa(\Add0~4_combout ),
	.datab(counter_reg_bit_0),
	.datac(\Add0~0_combout ),
	.datad(\Add0~2_combout ),
	.cin(gnd),
	.combout(\LessThan1~0_combout ),
	.cout());
defparam \LessThan1~0 .lut_mask = 16'hFFFE;
defparam \LessThan1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add0~6 (
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~5 ),
	.combout(\Add0~6_combout ),
	.cout(\Add0~7 ));
defparam \Add0~6 .lut_mask = 16'h5AAF;
defparam \Add0~6 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add0~8 (
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~7 ),
	.combout(\Add0~8_combout ),
	.cout(\Add0~9 ));
defparam \Add0~8 .lut_mask = 16'h5A5F;
defparam \Add0~8 .sum_lutc_input = "cin";

cycloneive_lcell_comb \LessThan1~1 (
	.dataa(\Add0~6_combout ),
	.datab(\Add0~8_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\LessThan1~1_combout ),
	.cout());
defparam \LessThan1~1 .lut_mask = 16'hEEEE;
defparam \LessThan1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add0~10 (
	.dataa(b_full),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~9 ),
	.combout(\Add0~10_combout ),
	.cout(\Add0~11 ));
defparam \Add0~10 .lut_mask = 16'h5AAF;
defparam \Add0~10 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add0~12 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add0~11 ),
	.combout(\Add0~12_combout ),
	.cout());
defparam \Add0~12 .lut_mask = 16'hF0F0;
defparam \Add0~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \LessThan1~2 (
	.dataa(\LessThan1~0_combout ),
	.datab(\LessThan1~1_combout ),
	.datac(\Add0~10_combout ),
	.datad(\Add0~12_combout ),
	.cin(gnd),
	.combout(\LessThan1~2_combout ),
	.cout());
defparam \LessThan1~2 .lut_mask = 16'h7FFF;
defparam \LessThan1~2 .sum_lutc_input = "datac";

dffeas fifo_AF(
	.clk(clk_clk),
	.d(\LessThan1~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_AF~q ),
	.prn(vcc));
defparam fifo_AF.is_wysiwyg = "true";
defparam fifo_AF.power_up = "low";

cycloneive_lcell_comb \ac~0 (
	.dataa(\nios_mcu_jtag_uart_0_alt_jtag_atlantic|t_ena~reg0_q ),
	.datab(\nios_mcu_jtag_uart_0_alt_jtag_atlantic|t_pause~reg0_q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ac~0_combout ),
	.cout());
defparam \ac~0 .lut_mask = 16'hEEEE;
defparam \ac~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ac~1 (
	.dataa(\ac~0_combout ),
	.datab(ac1),
	.datac(d_writedata_10),
	.datad(\ien_AE~0_combout ),
	.cin(gnd),
	.combout(\ac~1_combout ),
	.cout());
defparam \ac~1 .lut_mask = 16'hEFFF;
defparam \ac~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rvalid~0 (
	.dataa(b_non_empty),
	.datab(rvalid1),
	.datac(gnd),
	.datad(\fifo_rd~1_combout ),
	.cin(gnd),
	.combout(\rvalid~0_combout ),
	.cout());
defparam \rvalid~0 .lut_mask = 16'hAACC;
defparam \rvalid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \woverflow~0 (
	.dataa(rst1),
	.datab(m0_write),
	.datac(\av_waitrequest~0_combout ),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(\woverflow~0_combout ),
	.cout());
defparam \woverflow~0 .lut_mask = 16'hFEFF;
defparam \woverflow~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \woverflow~1 (
	.dataa(b_full1),
	.datab(woverflow1),
	.datac(gnd),
	.datad(\woverflow~0_combout ),
	.cin(gnd),
	.combout(\woverflow~1_combout ),
	.cout());
defparam \woverflow~1 .lut_mask = 16'hAACC;
defparam \woverflow~1 .sum_lutc_input = "datac";

endmodule

module nios_mcu_alt_jtag_atlantic (
	r_dat,
	adapted_tdo1,
	rst_n,
	rst11,
	t_dav,
	rvalid01,
	r_val,
	r_ena11,
	t_ena,
	wdata_0,
	t_pause,
	wdata_1,
	wdata_2,
	wdata_3,
	wdata_4,
	wdata_5,
	wdata_6,
	wdata_7,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	splitter_nodes_receive_0_3,
	virtual_ir_scan_reg,
	clr_reg,
	state_3,
	state_8,
	irf_reg_0_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	[7:0] r_dat;
output 	adapted_tdo1;
input 	rst_n;
output 	rst11;
input 	t_dav;
output 	rvalid01;
input 	r_val;
output 	r_ena11;
output 	t_ena;
output 	wdata_0;
output 	t_pause;
output 	wdata_1;
output 	wdata_2;
output 	wdata_3;
output 	wdata_4;
output 	wdata_5;
output 	wdata_6;
output 	wdata_7;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	splitter_nodes_receive_0_3;
input 	virtual_ir_scan_reg;
input 	clr_reg;
input 	state_3;
input 	state_8;
input 	irf_reg_0_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tck_t_dav~0_combout ;
wire \tck_t_dav~q ;
wire \state~1_combout ;
wire \always0~0_combout ;
wire \state~0_combout ;
wire \state~2_combout ;
wire \state~q ;
wire \count~9_combout ;
wire \td_shift[0]~4_combout ;
wire \count[2]~q ;
wire \count~8_combout ;
wire \count[3]~q ;
wire \count~7_combout ;
wire \count[4]~q ;
wire \count~6_combout ;
wire \count[5]~q ;
wire \count~5_combout ;
wire \count[6]~q ;
wire \count~4_combout ;
wire \count[7]~q ;
wire \count~2_combout ;
wire \count[8]~q ;
wire \count[9]~0_combout ;
wire \count[9]~q ;
wire \count~3_combout ;
wire \count[0]~q ;
wire \count~1_combout ;
wire \count[1]~q ;
wire \wdata[1]~2_combout ;
wire \user_saw_rvalid~0_combout ;
wire \user_saw_rvalid~q ;
wire \td_shift~10_combout ;
wire \td_shift[10]~q ;
wire \r_ena~0_combout ;
wire \rdata[7]~q ;
wire \td_shift~7_combout ;
wire \td_shift[9]~q ;
wire \td_shift~1_combout ;
wire \rdata[6]~q ;
wire \td_shift~21_combout ;
wire \td_shift[8]~q ;
wire \rdata[5]~q ;
wire \td_shift~19_combout ;
wire \td_shift~20_combout ;
wire \td_shift[7]~q ;
wire \rdata[4]~q ;
wire \td_shift~17_combout ;
wire \td_shift~18_combout ;
wire \td_shift[6]~q ;
wire \rdata[3]~q ;
wire \td_shift~15_combout ;
wire \td_shift~16_combout ;
wire \td_shift[5]~q ;
wire \rdata[2]~q ;
wire \td_shift~13_combout ;
wire \td_shift~14_combout ;
wire \td_shift[4]~q ;
wire \rdata[1]~q ;
wire \td_shift~11_combout ;
wire \td_shift~12_combout ;
wire \td_shift[3]~q ;
wire \rdata[0]~q ;
wire \td_shift~8_combout ;
wire \td_shift~9_combout ;
wire \td_shift[2]~q ;
wire \write_stalled~2_combout ;
wire \write_stalled~4_combout ;
wire \write_stalled~3_combout ;
wire \write_stalled~q ;
wire \td_shift~5_combout ;
wire \td_shift~6_combout ;
wire \td_shift[1]~q ;
wire \rvalid~q ;
wire \td_shift~0_combout ;
wire \td_shift~2_combout ;
wire \td_shift~3_combout ;
wire \td_shift[0]~q ;
wire \rvalid0~0_combout ;
wire \read~0_combout ;
wire \read~q ;
wire \read1~q ;
wire \read2~q ;
wire \read_req~q ;
wire \rvalid0~1_combout ;
wire \rst2~q ;
wire \rvalid0~2_combout ;
wire \write~0_combout ;
wire \wdata[1]~3_combout ;
wire \write~q ;
wire \write1~q ;
wire \write2~q ;
wire \write_valid~q ;
wire \t_ena~2_combout ;
wire \t_ena~3_combout ;
wire \always2~0_combout ;
wire \t_pause~0_combout ;
wire \jupdate~0_combout ;
wire \jupdate~q ;
wire \jupdate1~q ;
wire \jupdate2~q ;
wire \t_pause~1_combout ;


dffeas adapted_tdo(
	.clk(!altera_internal_jtag),
	.d(\td_shift[0]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(adapted_tdo1),
	.prn(vcc));
defparam adapted_tdo.is_wysiwyg = "true";
defparam adapted_tdo.power_up = "low";

dffeas rst1(
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rst11),
	.prn(vcc));
defparam rst1.is_wysiwyg = "true";
defparam rst1.power_up = "low";

dffeas rvalid0(
	.clk(clk),
	.d(\rvalid0~2_combout ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rvalid01),
	.prn(vcc));
defparam rvalid0.is_wysiwyg = "true";
defparam rvalid0.power_up = "low";

dffeas r_ena1(
	.clk(clk),
	.d(\rvalid0~0_combout ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_ena11),
	.prn(vcc));
defparam r_ena1.is_wysiwyg = "true";
defparam r_ena1.power_up = "low";

dffeas \t_ena~reg0 (
	.clk(clk),
	.d(\t_ena~3_combout ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(t_ena),
	.prn(vcc));
defparam \t_ena~reg0 .is_wysiwyg = "true";
defparam \t_ena~reg0 .power_up = "low";

dffeas \wdata[0] (
	.clk(altera_internal_jtag),
	.d(altera_internal_jtag1),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~3_combout ),
	.q(wdata_0),
	.prn(vcc));
defparam \wdata[0] .is_wysiwyg = "true";
defparam \wdata[0] .power_up = "low";

dffeas \t_pause~reg0 (
	.clk(clk),
	.d(\t_pause~1_combout ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(t_pause),
	.prn(vcc));
defparam \t_pause~reg0 .is_wysiwyg = "true";
defparam \t_pause~reg0 .power_up = "low";

dffeas \wdata[1] (
	.clk(altera_internal_jtag),
	.d(\td_shift[5]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~3_combout ),
	.q(wdata_1),
	.prn(vcc));
defparam \wdata[1] .is_wysiwyg = "true";
defparam \wdata[1] .power_up = "low";

dffeas \wdata[2] (
	.clk(altera_internal_jtag),
	.d(\td_shift[6]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~3_combout ),
	.q(wdata_2),
	.prn(vcc));
defparam \wdata[2] .is_wysiwyg = "true";
defparam \wdata[2] .power_up = "low";

dffeas \wdata[3] (
	.clk(altera_internal_jtag),
	.d(\td_shift[7]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~3_combout ),
	.q(wdata_3),
	.prn(vcc));
defparam \wdata[3] .is_wysiwyg = "true";
defparam \wdata[3] .power_up = "low";

dffeas \wdata[4] (
	.clk(altera_internal_jtag),
	.d(\td_shift[8]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~3_combout ),
	.q(wdata_4),
	.prn(vcc));
defparam \wdata[4] .is_wysiwyg = "true";
defparam \wdata[4] .power_up = "low";

dffeas \wdata[5] (
	.clk(altera_internal_jtag),
	.d(\td_shift[9]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~3_combout ),
	.q(wdata_5),
	.prn(vcc));
defparam \wdata[5] .is_wysiwyg = "true";
defparam \wdata[5] .power_up = "low";

dffeas \wdata[6] (
	.clk(altera_internal_jtag),
	.d(\td_shift[10]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~3_combout ),
	.q(wdata_6),
	.prn(vcc));
defparam \wdata[6] .is_wysiwyg = "true";
defparam \wdata[6] .power_up = "low";

dffeas \wdata[7] (
	.clk(altera_internal_jtag),
	.d(altera_internal_jtag1),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~3_combout ),
	.q(wdata_7),
	.prn(vcc));
defparam \wdata[7] .is_wysiwyg = "true";
defparam \wdata[7] .power_up = "low";

cycloneive_lcell_comb \tck_t_dav~0 (
	.dataa(t_dav),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\tck_t_dav~0_combout ),
	.cout());
defparam \tck_t_dav~0 .lut_mask = 16'h5555;
defparam \tck_t_dav~0 .sum_lutc_input = "datac";

dffeas tck_t_dav(
	.clk(altera_internal_jtag),
	.d(\tck_t_dav~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tck_t_dav~q ),
	.prn(vcc));
defparam tck_t_dav.is_wysiwyg = "true";
defparam tck_t_dav.power_up = "low";

cycloneive_lcell_comb \state~1 (
	.dataa(\state~q ),
	.datab(virtual_ir_scan_reg),
	.datac(splitter_nodes_receive_0_3),
	.datad(state_3),
	.cin(gnd),
	.combout(\state~1_combout ),
	.cout());
defparam \state~1 .lut_mask = 16'hEFFF;
defparam \state~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always0~0 (
	.dataa(splitter_nodes_receive_0_3),
	.datab(gnd),
	.datac(gnd),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\always0~0_combout ),
	.cout());
defparam \always0~0 .lut_mask = 16'hAAFF;
defparam \always0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \state~0 (
	.dataa(altera_internal_jtag1),
	.datab(gnd),
	.datac(irf_reg_0_1),
	.datad(\state~q ),
	.cin(gnd),
	.combout(\state~0_combout ),
	.cout());
defparam \state~0 .lut_mask = 16'hAFFF;
defparam \state~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \state~2 (
	.dataa(\state~1_combout ),
	.datab(state_4),
	.datac(\always0~0_combout ),
	.datad(\state~0_combout ),
	.cin(gnd),
	.combout(\state~2_combout ),
	.cout());
defparam \state~2 .lut_mask = 16'hFFFE;
defparam \state~2 .sum_lutc_input = "datac";

dffeas state(
	.clk(altera_internal_jtag),
	.d(\state~2_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state~q ),
	.prn(vcc));
defparam state.is_wysiwyg = "true";
defparam state.power_up = "low";

cycloneive_lcell_comb \count~9 (
	.dataa(\count[1]~q ),
	.datab(state_4),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~9_combout ),
	.cout());
defparam \count~9 .lut_mask = 16'hEEEE;
defparam \count~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift[0]~4 (
	.dataa(splitter_nodes_receive_0_3),
	.datab(state_4),
	.datac(state_3),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\td_shift[0]~4_combout ),
	.cout());
defparam \td_shift[0]~4 .lut_mask = 16'hFEFF;
defparam \td_shift[0]~4 .sum_lutc_input = "datac";

dffeas \count[2] (
	.clk(altera_internal_jtag),
	.d(\count~9_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[2]~q ),
	.prn(vcc));
defparam \count[2] .is_wysiwyg = "true";
defparam \count[2] .power_up = "low";

cycloneive_lcell_comb \count~8 (
	.dataa(state_4),
	.datab(\count[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~8_combout ),
	.cout());
defparam \count~8 .lut_mask = 16'hEEEE;
defparam \count~8 .sum_lutc_input = "datac";

dffeas \count[3] (
	.clk(altera_internal_jtag),
	.d(\count~8_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[3]~q ),
	.prn(vcc));
defparam \count[3] .is_wysiwyg = "true";
defparam \count[3] .power_up = "low";

cycloneive_lcell_comb \count~7 (
	.dataa(state_4),
	.datab(\count[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~7_combout ),
	.cout());
defparam \count~7 .lut_mask = 16'hEEEE;
defparam \count~7 .sum_lutc_input = "datac";

dffeas \count[4] (
	.clk(altera_internal_jtag),
	.d(\count~7_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[4]~q ),
	.prn(vcc));
defparam \count[4] .is_wysiwyg = "true";
defparam \count[4] .power_up = "low";

cycloneive_lcell_comb \count~6 (
	.dataa(state_4),
	.datab(\count[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~6_combout ),
	.cout());
defparam \count~6 .lut_mask = 16'hEEEE;
defparam \count~6 .sum_lutc_input = "datac";

dffeas \count[5] (
	.clk(altera_internal_jtag),
	.d(\count~6_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[5]~q ),
	.prn(vcc));
defparam \count[5] .is_wysiwyg = "true";
defparam \count[5] .power_up = "low";

cycloneive_lcell_comb \count~5 (
	.dataa(state_4),
	.datab(\count[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~5_combout ),
	.cout());
defparam \count~5 .lut_mask = 16'hEEEE;
defparam \count~5 .sum_lutc_input = "datac";

dffeas \count[6] (
	.clk(altera_internal_jtag),
	.d(\count~5_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[6]~q ),
	.prn(vcc));
defparam \count[6] .is_wysiwyg = "true";
defparam \count[6] .power_up = "low";

cycloneive_lcell_comb \count~4 (
	.dataa(state_4),
	.datab(\count[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~4_combout ),
	.cout());
defparam \count~4 .lut_mask = 16'hEEEE;
defparam \count~4 .sum_lutc_input = "datac";

dffeas \count[7] (
	.clk(altera_internal_jtag),
	.d(\count~4_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[7]~q ),
	.prn(vcc));
defparam \count[7] .is_wysiwyg = "true";
defparam \count[7] .power_up = "low";

cycloneive_lcell_comb \count~2 (
	.dataa(state_4),
	.datab(\count[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~2_combout ),
	.cout());
defparam \count~2 .lut_mask = 16'hEEEE;
defparam \count~2 .sum_lutc_input = "datac";

dffeas \count[8] (
	.clk(altera_internal_jtag),
	.d(\count~2_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[8]~q ),
	.prn(vcc));
defparam \count[8] .is_wysiwyg = "true";
defparam \count[8] .power_up = "low";

cycloneive_lcell_comb \count[9]~0 (
	.dataa(state_4),
	.datab(\state~0_combout ),
	.datac(\count[8]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\count[9]~0_combout ),
	.cout());
defparam \count[9]~0 .lut_mask = 16'h7F7F;
defparam \count[9]~0 .sum_lutc_input = "datac";

dffeas \count[9] (
	.clk(altera_internal_jtag),
	.d(\count[9]~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[9]~q ),
	.prn(vcc));
defparam \count[9] .is_wysiwyg = "true";
defparam \count[9] .power_up = "low";

cycloneive_lcell_comb \count~3 (
	.dataa(state_4),
	.datab(gnd),
	.datac(gnd),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\count~3_combout ),
	.cout());
defparam \count~3 .lut_mask = 16'hAAFF;
defparam \count~3 .sum_lutc_input = "datac";

dffeas \count[0] (
	.clk(altera_internal_jtag),
	.d(\count~3_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[0]~q ),
	.prn(vcc));
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";

cycloneive_lcell_comb \count~1 (
	.dataa(state_4),
	.datab(\count[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~1_combout ),
	.cout());
defparam \count~1 .lut_mask = 16'hEEEE;
defparam \count~1 .sum_lutc_input = "datac";

dffeas \count[1] (
	.clk(altera_internal_jtag),
	.d(\count~1_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\count[1]~q ),
	.prn(vcc));
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";

cycloneive_lcell_comb \wdata[1]~2 (
	.dataa(\state~q ),
	.datab(state_4),
	.datac(\always0~0_combout ),
	.datad(irf_reg_0_1),
	.cin(gnd),
	.combout(\wdata[1]~2_combout ),
	.cout());
defparam \wdata[1]~2 .lut_mask = 16'hFEFF;
defparam \wdata[1]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \user_saw_rvalid~0 (
	.dataa(\td_shift[0]~q ),
	.datab(\user_saw_rvalid~q ),
	.datac(\count[0]~q ),
	.datad(\wdata[1]~2_combout ),
	.cin(gnd),
	.combout(\user_saw_rvalid~0_combout ),
	.cout());
defparam \user_saw_rvalid~0 .lut_mask = 16'hEFFE;
defparam \user_saw_rvalid~0 .sum_lutc_input = "datac";

dffeas user_saw_rvalid(
	.clk(altera_internal_jtag),
	.d(\user_saw_rvalid~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\user_saw_rvalid~q ),
	.prn(vcc));
defparam user_saw_rvalid.is_wysiwyg = "true";
defparam user_saw_rvalid.power_up = "low";

cycloneive_lcell_comb \td_shift~10 (
	.dataa(altera_internal_jtag1),
	.datab(state_4),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\td_shift~10_combout ),
	.cout());
defparam \td_shift~10 .lut_mask = 16'hEEEE;
defparam \td_shift~10 .sum_lutc_input = "datac";

dffeas \td_shift[10] (
	.clk(altera_internal_jtag),
	.d(\td_shift~10_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[10]~q ),
	.prn(vcc));
defparam \td_shift[10] .is_wysiwyg = "true";
defparam \td_shift[10] .power_up = "low";

cycloneive_lcell_comb \r_ena~0 (
	.dataa(r_val),
	.datab(r_ena11),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\r_ena~0_combout ),
	.cout());
defparam \r_ena~0 .lut_mask = 16'hEEEE;
defparam \r_ena~0 .sum_lutc_input = "datac";

dffeas \rdata[7] (
	.clk(clk),
	.d(r_dat[7]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[7]~q ),
	.prn(vcc));
defparam \rdata[7] .is_wysiwyg = "true";
defparam \rdata[7] .power_up = "low";

cycloneive_lcell_comb \td_shift~7 (
	.dataa(\td_shift[10]~q ),
	.datab(\rdata[7]~q ),
	.datac(gnd),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\td_shift~7_combout ),
	.cout());
defparam \td_shift~7 .lut_mask = 16'hAACC;
defparam \td_shift~7 .sum_lutc_input = "datac";

dffeas \td_shift[9] (
	.clk(altera_internal_jtag),
	.d(\td_shift~7_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[9]~q ),
	.prn(vcc));
defparam \td_shift[9] .is_wysiwyg = "true";
defparam \td_shift[9] .power_up = "low";

cycloneive_lcell_comb \td_shift~1 (
	.dataa(\state~q ),
	.datab(\count[1]~q ),
	.datac(\user_saw_rvalid~q ),
	.datad(\td_shift[9]~q ),
	.cin(gnd),
	.combout(\td_shift~1_combout ),
	.cout());
defparam \td_shift~1 .lut_mask = 16'hEFFF;
defparam \td_shift~1 .sum_lutc_input = "datac";

dffeas \rdata[6] (
	.clk(clk),
	.d(r_dat[6]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[6]~q ),
	.prn(vcc));
defparam \rdata[6] .is_wysiwyg = "true";
defparam \rdata[6] .power_up = "low";

cycloneive_lcell_comb \td_shift~21 (
	.dataa(\td_shift[9]~q ),
	.datab(\rdata[6]~q ),
	.datac(gnd),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\td_shift~21_combout ),
	.cout());
defparam \td_shift~21 .lut_mask = 16'hAACC;
defparam \td_shift~21 .sum_lutc_input = "datac";

dffeas \td_shift[8] (
	.clk(altera_internal_jtag),
	.d(\td_shift~21_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[8]~q ),
	.prn(vcc));
defparam \td_shift[8] .is_wysiwyg = "true";
defparam \td_shift[8] .power_up = "low";

dffeas \rdata[5] (
	.clk(clk),
	.d(r_dat[5]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[5]~q ),
	.prn(vcc));
defparam \rdata[5] .is_wysiwyg = "true";
defparam \rdata[5] .power_up = "low";

cycloneive_lcell_comb \td_shift~19 (
	.dataa(\td_shift[8]~q ),
	.datab(\rdata[5]~q ),
	.datac(\count[9]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\td_shift~19_combout ),
	.cout());
defparam \td_shift~19 .lut_mask = 16'hACAC;
defparam \td_shift~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift~20 (
	.dataa(state_4),
	.datab(irf_reg_0_1),
	.datac(\td_shift~1_combout ),
	.datad(\td_shift~19_combout ),
	.cin(gnd),
	.combout(\td_shift~20_combout ),
	.cout());
defparam \td_shift~20 .lut_mask = 16'hFFEF;
defparam \td_shift~20 .sum_lutc_input = "datac";

dffeas \td_shift[7] (
	.clk(altera_internal_jtag),
	.d(\td_shift~20_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[7]~q ),
	.prn(vcc));
defparam \td_shift[7] .is_wysiwyg = "true";
defparam \td_shift[7] .power_up = "low";

dffeas \rdata[4] (
	.clk(clk),
	.d(r_dat[4]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[4]~q ),
	.prn(vcc));
defparam \rdata[4] .is_wysiwyg = "true";
defparam \rdata[4] .power_up = "low";

cycloneive_lcell_comb \td_shift~17 (
	.dataa(\td_shift[7]~q ),
	.datab(\rdata[4]~q ),
	.datac(gnd),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\td_shift~17_combout ),
	.cout());
defparam \td_shift~17 .lut_mask = 16'hAACC;
defparam \td_shift~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift~18 (
	.dataa(irf_reg_0_1),
	.datab(\td_shift~17_combout ),
	.datac(state_4),
	.datad(\td_shift~1_combout ),
	.cin(gnd),
	.combout(\td_shift~18_combout ),
	.cout());
defparam \td_shift~18 .lut_mask = 16'hACFF;
defparam \td_shift~18 .sum_lutc_input = "datac";

dffeas \td_shift[6] (
	.clk(altera_internal_jtag),
	.d(\td_shift~18_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[6]~q ),
	.prn(vcc));
defparam \td_shift[6] .is_wysiwyg = "true";
defparam \td_shift[6] .power_up = "low";

dffeas \rdata[3] (
	.clk(clk),
	.d(r_dat[3]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[3]~q ),
	.prn(vcc));
defparam \rdata[3] .is_wysiwyg = "true";
defparam \rdata[3] .power_up = "low";

cycloneive_lcell_comb \td_shift~15 (
	.dataa(\td_shift[6]~q ),
	.datab(\rdata[3]~q ),
	.datac(gnd),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\td_shift~15_combout ),
	.cout());
defparam \td_shift~15 .lut_mask = 16'hAACC;
defparam \td_shift~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift~16 (
	.dataa(irf_reg_0_1),
	.datab(\td_shift~15_combout ),
	.datac(state_4),
	.datad(\td_shift~1_combout ),
	.cin(gnd),
	.combout(\td_shift~16_combout ),
	.cout());
defparam \td_shift~16 .lut_mask = 16'hACFF;
defparam \td_shift~16 .sum_lutc_input = "datac";

dffeas \td_shift[5] (
	.clk(altera_internal_jtag),
	.d(\td_shift~16_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[5]~q ),
	.prn(vcc));
defparam \td_shift[5] .is_wysiwyg = "true";
defparam \td_shift[5] .power_up = "low";

dffeas \rdata[2] (
	.clk(clk),
	.d(r_dat[2]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[2]~q ),
	.prn(vcc));
defparam \rdata[2] .is_wysiwyg = "true";
defparam \rdata[2] .power_up = "low";

cycloneive_lcell_comb \td_shift~13 (
	.dataa(\td_shift[5]~q ),
	.datab(\rdata[2]~q ),
	.datac(\count[9]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\td_shift~13_combout ),
	.cout());
defparam \td_shift~13 .lut_mask = 16'hACAC;
defparam \td_shift~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift~14 (
	.dataa(state_4),
	.datab(irf_reg_0_1),
	.datac(\td_shift~1_combout ),
	.datad(\td_shift~13_combout ),
	.cin(gnd),
	.combout(\td_shift~14_combout ),
	.cout());
defparam \td_shift~14 .lut_mask = 16'hFFEF;
defparam \td_shift~14 .sum_lutc_input = "datac";

dffeas \td_shift[4] (
	.clk(altera_internal_jtag),
	.d(\td_shift~14_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[4]~q ),
	.prn(vcc));
defparam \td_shift[4] .is_wysiwyg = "true";
defparam \td_shift[4] .power_up = "low";

dffeas \rdata[1] (
	.clk(clk),
	.d(r_dat[1]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[1]~q ),
	.prn(vcc));
defparam \rdata[1] .is_wysiwyg = "true";
defparam \rdata[1] .power_up = "low";

cycloneive_lcell_comb \td_shift~11 (
	.dataa(\td_shift[4]~q ),
	.datab(\rdata[1]~q ),
	.datac(\count[9]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\td_shift~11_combout ),
	.cout());
defparam \td_shift~11 .lut_mask = 16'hACAC;
defparam \td_shift~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift~12 (
	.dataa(state_4),
	.datab(irf_reg_0_1),
	.datac(\td_shift~1_combout ),
	.datad(\td_shift~11_combout ),
	.cin(gnd),
	.combout(\td_shift~12_combout ),
	.cout());
defparam \td_shift~12 .lut_mask = 16'hFFEF;
defparam \td_shift~12 .sum_lutc_input = "datac";

dffeas \td_shift[3] (
	.clk(altera_internal_jtag),
	.d(\td_shift~12_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[3]~q ),
	.prn(vcc));
defparam \td_shift[3] .is_wysiwyg = "true";
defparam \td_shift[3] .power_up = "low";

dffeas \rdata[0] (
	.clk(clk),
	.d(r_dat[0]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[0]~q ),
	.prn(vcc));
defparam \rdata[0] .is_wysiwyg = "true";
defparam \rdata[0] .power_up = "low";

cycloneive_lcell_comb \td_shift~8 (
	.dataa(\td_shift[3]~q ),
	.datab(\rdata[0]~q ),
	.datac(gnd),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\td_shift~8_combout ),
	.cout());
defparam \td_shift~8 .lut_mask = 16'hAACC;
defparam \td_shift~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift~9 (
	.dataa(irf_reg_0_1),
	.datab(\td_shift~8_combout ),
	.datac(state_4),
	.datad(\td_shift~1_combout ),
	.cin(gnd),
	.combout(\td_shift~9_combout ),
	.cout());
defparam \td_shift~9 .lut_mask = 16'hACFF;
defparam \td_shift~9 .sum_lutc_input = "datac";

dffeas \td_shift[2] (
	.clk(altera_internal_jtag),
	.d(\td_shift~9_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[2]~q ),
	.prn(vcc));
defparam \td_shift[2] .is_wysiwyg = "true";
defparam \td_shift[2] .power_up = "low";

cycloneive_lcell_comb \write_stalled~2 (
	.dataa(\write_stalled~q ),
	.datab(\td_shift[10]~q ),
	.datac(altera_internal_jtag1),
	.datad(\tck_t_dav~q ),
	.cin(gnd),
	.combout(\write_stalled~2_combout ),
	.cout());
defparam \write_stalled~2 .lut_mask = 16'hEFFF;
defparam \write_stalled~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \write_stalled~4 (
	.dataa(splitter_nodes_receive_0_3),
	.datab(virtual_ir_scan_reg),
	.datac(irf_reg_0_1),
	.datad(gnd),
	.cin(gnd),
	.combout(\write_stalled~4_combout ),
	.cout());
defparam \write_stalled~4 .lut_mask = 16'hBFBF;
defparam \write_stalled~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \write_stalled~3 (
	.dataa(\count[1]~q ),
	.datab(\state~q ),
	.datac(state_4),
	.datad(\write_stalled~4_combout ),
	.cin(gnd),
	.combout(\write_stalled~3_combout ),
	.cout());
defparam \write_stalled~3 .lut_mask = 16'hFFFE;
defparam \write_stalled~3 .sum_lutc_input = "datac";

dffeas write_stalled(
	.clk(altera_internal_jtag),
	.d(\write_stalled~2_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~3_combout ),
	.q(\write_stalled~q ),
	.prn(vcc));
defparam write_stalled.is_wysiwyg = "true";
defparam write_stalled.power_up = "low";

cycloneive_lcell_comb \td_shift~5 (
	.dataa(\td_shift[2]~q ),
	.datab(\write_stalled~q ),
	.datac(gnd),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\td_shift~5_combout ),
	.cout());
defparam \td_shift~5 .lut_mask = 16'hAACC;
defparam \td_shift~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift~6 (
	.dataa(irf_reg_0_1),
	.datab(\td_shift~5_combout ),
	.datac(state_4),
	.datad(\td_shift~1_combout ),
	.cin(gnd),
	.combout(\td_shift~6_combout ),
	.cout());
defparam \td_shift~6 .lut_mask = 16'hACFF;
defparam \td_shift~6 .sum_lutc_input = "datac";

dffeas \td_shift[1] (
	.clk(altera_internal_jtag),
	.d(\td_shift~6_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[1]~q ),
	.prn(vcc));
defparam \td_shift[1] .is_wysiwyg = "true";
defparam \td_shift[1] .power_up = "low";

dffeas rvalid(
	.clk(clk),
	.d(rvalid01),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rvalid~q ),
	.prn(vcc));
defparam rvalid.is_wysiwyg = "true";
defparam rvalid.power_up = "low";

cycloneive_lcell_comb \td_shift~0 (
	.dataa(\td_shift[1]~q ),
	.datab(\rvalid~q ),
	.datac(gnd),
	.datad(\count[9]~q ),
	.cin(gnd),
	.combout(\td_shift~0_combout ),
	.cout());
defparam \td_shift~0 .lut_mask = 16'hAACC;
defparam \td_shift~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift~2 (
	.dataa(\td_shift~1_combout ),
	.datab(altera_internal_jtag1),
	.datac(\state~q ),
	.datad(irf_reg_0_1),
	.cin(gnd),
	.combout(\td_shift~2_combout ),
	.cout());
defparam \td_shift~2 .lut_mask = 16'hEFFF;
defparam \td_shift~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \td_shift~3 (
	.dataa(\tck_t_dav~q ),
	.datab(\td_shift~0_combout ),
	.datac(\td_shift~2_combout ),
	.datad(\state~q ),
	.cin(gnd),
	.combout(\td_shift~3_combout ),
	.cout());
defparam \td_shift~3 .lut_mask = 16'hACFF;
defparam \td_shift~3 .sum_lutc_input = "datac";

dffeas \td_shift[0] (
	.clk(altera_internal_jtag),
	.d(\td_shift~3_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~4_combout ),
	.q(\td_shift[0]~q ),
	.prn(vcc));
defparam \td_shift[0] .is_wysiwyg = "true";
defparam \td_shift[0] .power_up = "low";

cycloneive_lcell_comb \rvalid0~0 (
	.dataa(rvalid01),
	.datab(r_val),
	.datac(r_ena11),
	.datad(gnd),
	.cin(gnd),
	.combout(\rvalid0~0_combout ),
	.cout());
defparam \rvalid0~0 .lut_mask = 16'h7F7F;
defparam \rvalid0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read~0 (
	.dataa(\read~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\read~0_combout ),
	.cout());
defparam \read~0 .lut_mask = 16'h5555;
defparam \read~0 .sum_lutc_input = "datac";

dffeas read(
	.clk(altera_internal_jtag),
	.d(\read~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~3_combout ),
	.q(\read~q ),
	.prn(vcc));
defparam read.is_wysiwyg = "true";
defparam read.power_up = "low";

dffeas read1(
	.clk(clk),
	.d(\read~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read1~q ),
	.prn(vcc));
defparam read1.is_wysiwyg = "true";
defparam read1.power_up = "low";

dffeas read2(
	.clk(clk),
	.d(\read1~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read2~q ),
	.prn(vcc));
defparam read2.is_wysiwyg = "true";
defparam read2.power_up = "low";

dffeas read_req(
	.clk(altera_internal_jtag),
	.d(\td_shift[9]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~3_combout ),
	.q(\read_req~q ),
	.prn(vcc));
defparam read_req.is_wysiwyg = "true";
defparam read_req.power_up = "low";

cycloneive_lcell_comb \rvalid0~1 (
	.dataa(\read1~q ),
	.datab(\read2~q ),
	.datac(\user_saw_rvalid~q ),
	.datad(\read_req~q ),
	.cin(gnd),
	.combout(\rvalid0~1_combout ),
	.cout());
defparam \rvalid0~1 .lut_mask = 16'h6FFF;
defparam \rvalid0~1 .sum_lutc_input = "datac";

dffeas rst2(
	.clk(clk),
	.d(rst11),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rst2~q ),
	.prn(vcc));
defparam rst2.is_wysiwyg = "true";
defparam rst2.power_up = "low";

cycloneive_lcell_comb \rvalid0~2 (
	.dataa(\rvalid0~0_combout ),
	.datab(\rvalid0~1_combout ),
	.datac(gnd),
	.datad(\rst2~q ),
	.cin(gnd),
	.combout(\rvalid0~2_combout ),
	.cout());
defparam \rvalid0~2 .lut_mask = 16'hDDFF;
defparam \rvalid0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \write~0 (
	.dataa(\write~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\write~0_combout ),
	.cout());
defparam \write~0 .lut_mask = 16'h5555;
defparam \write~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wdata[1]~3 (
	.dataa(\count[8]~q ),
	.datab(\state~q ),
	.datac(state_4),
	.datad(\write_stalled~4_combout ),
	.cin(gnd),
	.combout(\wdata[1]~3_combout ),
	.cout());
defparam \wdata[1]~3 .lut_mask = 16'hFFFE;
defparam \wdata[1]~3 .sum_lutc_input = "datac";

dffeas write(
	.clk(altera_internal_jtag),
	.d(\write~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[1]~3_combout ),
	.q(\write~q ),
	.prn(vcc));
defparam write.is_wysiwyg = "true";
defparam write.power_up = "low";

dffeas write1(
	.clk(clk),
	.d(\write~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\write1~q ),
	.prn(vcc));
defparam write1.is_wysiwyg = "true";
defparam write1.power_up = "low";

dffeas write2(
	.clk(clk),
	.d(\write1~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\write2~q ),
	.prn(vcc));
defparam write2.is_wysiwyg = "true";
defparam write2.power_up = "low";

dffeas write_valid(
	.clk(altera_internal_jtag),
	.d(\td_shift[10]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~3_combout ),
	.q(\write_valid~q ),
	.prn(vcc));
defparam write_valid.is_wysiwyg = "true";
defparam write_valid.power_up = "low";

cycloneive_lcell_comb \t_ena~2 (
	.dataa(t_ena),
	.datab(\write_valid~q ),
	.datac(t_dav),
	.datad(\write_stalled~q ),
	.cin(gnd),
	.combout(\t_ena~2_combout ),
	.cout());
defparam \t_ena~2 .lut_mask = 16'hEFFF;
defparam \t_ena~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \t_ena~3 (
	.dataa(\write1~q ),
	.datab(\write2~q ),
	.datac(\rst2~q ),
	.datad(\t_ena~2_combout ),
	.cin(gnd),
	.combout(\t_ena~3_combout ),
	.cout());
defparam \t_ena~3 .lut_mask = 16'hFFF6;
defparam \t_ena~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always2~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\write1~q ),
	.datad(\write2~q ),
	.cin(gnd),
	.combout(\always2~0_combout ),
	.cout());
defparam \always2~0 .lut_mask = 16'h0FF0;
defparam \always2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \t_pause~0 (
	.dataa(\always2~0_combout ),
	.datab(t_dav),
	.datac(\write_stalled~q ),
	.datad(\write_valid~q ),
	.cin(gnd),
	.combout(\t_pause~0_combout ),
	.cout());
defparam \t_pause~0 .lut_mask = 16'hFEFF;
defparam \t_pause~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \jupdate~0 (
	.dataa(\jupdate~q ),
	.datab(irf_reg_0_1),
	.datac(\always0~0_combout ),
	.datad(state_8),
	.cin(gnd),
	.combout(\jupdate~0_combout ),
	.cout());
defparam \jupdate~0 .lut_mask = 16'h6996;
defparam \jupdate~0 .sum_lutc_input = "datac";

dffeas jupdate(
	.clk(!altera_internal_jtag),
	.d(\jupdate~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jupdate~q ),
	.prn(vcc));
defparam jupdate.is_wysiwyg = "true";
defparam jupdate.power_up = "low";

dffeas jupdate1(
	.clk(clk),
	.d(\jupdate~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jupdate1~q ),
	.prn(vcc));
defparam jupdate1.is_wysiwyg = "true";
defparam jupdate1.power_up = "low";

dffeas jupdate2(
	.clk(clk),
	.d(\jupdate1~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jupdate2~q ),
	.prn(vcc));
defparam jupdate2.is_wysiwyg = "true";
defparam jupdate2.power_up = "low";

cycloneive_lcell_comb \t_pause~1 (
	.dataa(\rst2~q ),
	.datab(\t_pause~0_combout ),
	.datac(\jupdate1~q ),
	.datad(\jupdate2~q ),
	.cin(gnd),
	.combout(\t_pause~1_combout ),
	.cout());
defparam \t_pause~1 .lut_mask = 16'hEFFE;
defparam \t_pause~1 .sum_lutc_input = "datac";

endmodule

module nios_mcu_nios_mcu_jtag_uart_0_scfifo_r (
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	r_sync_rst,
	b_full,
	b_non_empty,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	t_ena,
	fifo_rd,
	wr_rfifo,
	wdata_0,
	fifo_rd1,
	wdata_1,
	wdata_2,
	wdata_3,
	wdata_4,
	wdata_5,
	wdata_6,
	wdata_7,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
input 	r_sync_rst;
output 	b_full;
output 	b_non_empty;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	t_ena;
input 	fifo_rd;
input 	wr_rfifo;
input 	wdata_0;
input 	fifo_rd1;
input 	wdata_1;
input 	wdata_2;
input 	wdata_3;
input 	wdata_4;
input 	wdata_5;
input 	wdata_6;
input 	wdata_7;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nios_mcu_scfifo_1 rfifo(
	.q({q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.r_sync_rst(r_sync_rst),
	.b_full(b_full),
	.b_non_empty(b_non_empty),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.t_ena(t_ena),
	.fifo_rd(fifo_rd),
	.wrreq(wr_rfifo),
	.data({wdata_7,wdata_6,wdata_5,wdata_4,wdata_3,wdata_2,wdata_1,wdata_0}),
	.fifo_rd1(fifo_rd1),
	.clock(clk_clk));

endmodule

module nios_mcu_scfifo_1 (
	q,
	r_sync_rst,
	b_full,
	b_non_empty,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	t_ena,
	fifo_rd,
	wrreq,
	data,
	fifo_rd1,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	r_sync_rst;
output 	b_full;
output 	b_non_empty;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	t_ena;
input 	fifo_rd;
input 	wrreq;
input 	[7:0] data;
input 	fifo_rd1;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nios_mcu_scfifo_jr21 auto_generated(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.r_sync_rst(r_sync_rst),
	.b_full(b_full),
	.b_non_empty(b_non_empty),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.t_ena(t_ena),
	.fifo_rd(fifo_rd),
	.wrreq(wrreq),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.fifo_rd1(fifo_rd1),
	.clock(clock));

endmodule

module nios_mcu_scfifo_jr21 (
	q,
	r_sync_rst,
	b_full,
	b_non_empty,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	t_ena,
	fifo_rd,
	wrreq,
	data,
	fifo_rd1,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	r_sync_rst;
output 	b_full;
output 	b_non_empty;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	t_ena;
input 	fifo_rd;
input 	wrreq;
input 	[7:0] data;
input 	fifo_rd1;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nios_mcu_a_dpfifo_l011 dpfifo(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.r_sync_rst(r_sync_rst),
	.b_full(b_full),
	.b_non_empty(b_non_empty),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.t_ena(t_ena),
	.fifo_rd(fifo_rd),
	.wreq(wrreq),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.fifo_rd1(fifo_rd1),
	.clock(clock));

endmodule

module nios_mcu_a_dpfifo_l011 (
	q,
	r_sync_rst,
	b_full,
	b_non_empty,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	t_ena,
	fifo_rd,
	wreq,
	data,
	fifo_rd1,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	r_sync_rst;
output 	b_full;
output 	b_non_empty;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	t_ena;
input 	fifo_rd;
input 	wreq;
input 	[7:0] data;
input 	fifo_rd1;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \wr_ptr|counter_reg_bit[5]~q ;
wire \rd_ptr_count|counter_reg_bit[0]~q ;
wire \rd_ptr_count|counter_reg_bit[1]~q ;
wire \rd_ptr_count|counter_reg_bit[2]~q ;
wire \rd_ptr_count|counter_reg_bit[3]~q ;
wire \rd_ptr_count|counter_reg_bit[4]~q ;
wire \rd_ptr_count|counter_reg_bit[5]~q ;


nios_mcu_cntr_1ob_1 wr_ptr(
	.r_sync_rst(r_sync_rst),
	.wr_rfifo(wreq),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\wr_ptr|counter_reg_bit[5]~q ),
	.clock(clock));

nios_mcu_cntr_1ob rd_ptr_count(
	.r_sync_rst(r_sync_rst),
	.fifo_rd(fifo_rd),
	.counter_reg_bit_0(\rd_ptr_count|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_count|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_count|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_count|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\rd_ptr_count|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\rd_ptr_count|counter_reg_bit[5]~q ),
	.clock(clock));

nios_mcu_altsyncram_nio1 FIFOram(
	.q_b({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.clocken1(fifo_rd),
	.wren_a(wreq),
	.data_a({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.address_a({\wr_ptr|counter_reg_bit[5]~q ,\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.address_b({\rd_ptr_count|counter_reg_bit[5]~q ,\rd_ptr_count|counter_reg_bit[4]~q ,\rd_ptr_count|counter_reg_bit[3]~q ,\rd_ptr_count|counter_reg_bit[2]~q ,\rd_ptr_count|counter_reg_bit[1]~q ,\rd_ptr_count|counter_reg_bit[0]~q }),
	.clock0(clock),
	.clock1(clock));

nios_mcu_a_fefifo_7cf fifo_state(
	.r_sync_rst(r_sync_rst),
	.b_full1(b_full),
	.b_non_empty1(b_non_empty),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.t_ena(t_ena),
	.fifo_rd(fifo_rd),
	.wreq(wreq),
	.fifo_rd1(fifo_rd1),
	.clock(clock));

endmodule

module nios_mcu_a_fefifo_7cf (
	r_sync_rst,
	b_full1,
	b_non_empty1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	t_ena,
	fifo_rd,
	wreq,
	fifo_rd1,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
output 	b_full1;
output 	b_non_empty1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	t_ena;
input 	fifo_rd;
input 	wreq;
input 	fifo_rd1;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \_~4_combout ;
wire \b_full~0_combout ;
wire \b_full~1_combout ;
wire \b_full~2_combout ;
wire \b_non_empty~0_combout ;
wire \_~2_combout ;
wire \_~3_combout ;
wire \b_non_empty~1_combout ;


nios_mcu_cntr_do7 count_usedw(
	.r_sync_rst(r_sync_rst),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.updown(wreq),
	._(\_~4_combout ),
	.clock(clock));

cycloneive_lcell_comb \_~4 (
	.dataa(t_ena),
	.datab(b_full1),
	.datac(b_non_empty1),
	.datad(fifo_rd1),
	.cin(gnd),
	.combout(\_~4_combout ),
	.cout());
defparam \_~4 .lut_mask = 16'h6996;
defparam \_~4 .sum_lutc_input = "datac";

dffeas b_full(
	.clk(clock),
	.d(\b_full~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_full1),
	.prn(vcc));
defparam b_full.is_wysiwyg = "true";
defparam b_full.power_up = "low";

dffeas b_non_empty(
	.clk(clock),
	.d(\b_non_empty~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_non_empty1),
	.prn(vcc));
defparam b_non_empty.is_wysiwyg = "true";
defparam b_non_empty.power_up = "low";

cycloneive_lcell_comb \b_full~0 (
	.dataa(b_non_empty1),
	.datab(counter_reg_bit_5),
	.datac(counter_reg_bit_4),
	.datad(counter_reg_bit_3),
	.cin(gnd),
	.combout(\b_full~0_combout ),
	.cout());
defparam \b_full~0 .lut_mask = 16'hFFFE;
defparam \b_full~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_full~1 (
	.dataa(counter_reg_bit_2),
	.datab(counter_reg_bit_1),
	.datac(counter_reg_bit_0),
	.datad(t_ena),
	.cin(gnd),
	.combout(\b_full~1_combout ),
	.cout());
defparam \b_full~1 .lut_mask = 16'hFFFE;
defparam \b_full~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_full~2 (
	.dataa(b_full1),
	.datab(\b_full~0_combout ),
	.datac(\b_full~1_combout ),
	.datad(fifo_rd),
	.cin(gnd),
	.combout(\b_full~2_combout ),
	.cout());
defparam \b_full~2 .lut_mask = 16'hFEFF;
defparam \b_full~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_non_empty~0 (
	.dataa(b_full1),
	.datab(t_ena),
	.datac(gnd),
	.datad(b_non_empty1),
	.cin(gnd),
	.combout(\b_non_empty~0_combout ),
	.cout());
defparam \b_non_empty~0 .lut_mask = 16'hEEFF;
defparam \b_non_empty~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~2 (
	.dataa(counter_reg_bit_3),
	.datab(counter_reg_bit_2),
	.datac(counter_reg_bit_1),
	.datad(counter_reg_bit_0),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hFEFF;
defparam \_~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~3 (
	.dataa(counter_reg_bit_5),
	.datab(counter_reg_bit_4),
	.datac(wreq),
	.datad(\_~2_combout ),
	.cin(gnd),
	.combout(\_~3_combout ),
	.cout());
defparam \_~3 .lut_mask = 16'hFFFE;
defparam \_~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_non_empty~1 (
	.dataa(\b_non_empty~0_combout ),
	.datab(b_non_empty1),
	.datac(\_~3_combout ),
	.datad(fifo_rd1),
	.cin(gnd),
	.combout(\b_non_empty~1_combout ),
	.cout());
defparam \b_non_empty~1 .lut_mask = 16'hFEFF;
defparam \b_non_empty~1 .sum_lutc_input = "datac";

endmodule

module nios_mcu_cntr_do7 (
	r_sync_rst,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	updown,
	_,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	updown;
input 	_;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita0~combout ;


dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A6F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5A6F;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout());
defparam counter_comb_bita5.lut_mask = 16'h5A5A;
defparam counter_comb_bita5.sum_lutc_input = "cin";

endmodule

module nios_mcu_altsyncram_nio1 (
	q_b,
	clocken1,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock0,
	clock1)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q_b;
input 	clocken1;
input 	wren_a;
input 	[7:0] data_a;
input 	[5:0] address_a;
input 	[5:0] address_b;
input 	clock0;
input 	clock1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk1_core_clock_enable = "ena1";
defparam ram_block1a0.clk1_input_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "nios_mcu_jtag_uart_0:jtag_uart_0|nios_mcu_jtag_uart_0_scfifo_r:the_nios_mcu_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_jr21:auto_generated|a_dpfifo_l011:dpfifo|altsyncram_nio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 6;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 63;
defparam ram_block1a0.port_a_logical_ram_depth = 64;
defparam ram_block1a0.port_a_logical_ram_width = 8;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 6;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 63;
defparam ram_block1a0.port_b_logical_ram_depth = 64;
defparam ram_block1a0.port_b_logical_ram_width = 8;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cycloneive_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk1_core_clock_enable = "ena1";
defparam ram_block1a1.clk1_input_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "nios_mcu_jtag_uart_0:jtag_uart_0|nios_mcu_jtag_uart_0_scfifo_r:the_nios_mcu_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_jr21:auto_generated|a_dpfifo_l011:dpfifo|altsyncram_nio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 6;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 63;
defparam ram_block1a1.port_a_logical_ram_depth = 64;
defparam ram_block1a1.port_a_logical_ram_width = 8;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 6;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 63;
defparam ram_block1a1.port_b_logical_ram_depth = 64;
defparam ram_block1a1.port_b_logical_ram_width = 8;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cycloneive_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk1_core_clock_enable = "ena1";
defparam ram_block1a2.clk1_input_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "nios_mcu_jtag_uart_0:jtag_uart_0|nios_mcu_jtag_uart_0_scfifo_r:the_nios_mcu_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_jr21:auto_generated|a_dpfifo_l011:dpfifo|altsyncram_nio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 6;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 63;
defparam ram_block1a2.port_a_logical_ram_depth = 64;
defparam ram_block1a2.port_a_logical_ram_width = 8;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 6;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 63;
defparam ram_block1a2.port_b_logical_ram_depth = 64;
defparam ram_block1a2.port_b_logical_ram_width = 8;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cycloneive_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk1_core_clock_enable = "ena1";
defparam ram_block1a3.clk1_input_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "nios_mcu_jtag_uart_0:jtag_uart_0|nios_mcu_jtag_uart_0_scfifo_r:the_nios_mcu_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_jr21:auto_generated|a_dpfifo_l011:dpfifo|altsyncram_nio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 6;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 63;
defparam ram_block1a3.port_a_logical_ram_depth = 64;
defparam ram_block1a3.port_a_logical_ram_width = 8;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 6;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 63;
defparam ram_block1a3.port_b_logical_ram_depth = 64;
defparam ram_block1a3.port_b_logical_ram_width = 8;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cycloneive_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk1_core_clock_enable = "ena1";
defparam ram_block1a4.clk1_input_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "nios_mcu_jtag_uart_0:jtag_uart_0|nios_mcu_jtag_uart_0_scfifo_r:the_nios_mcu_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_jr21:auto_generated|a_dpfifo_l011:dpfifo|altsyncram_nio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 6;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 63;
defparam ram_block1a4.port_a_logical_ram_depth = 64;
defparam ram_block1a4.port_a_logical_ram_width = 8;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 6;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 63;
defparam ram_block1a4.port_b_logical_ram_depth = 64;
defparam ram_block1a4.port_b_logical_ram_width = 8;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk1_core_clock_enable = "ena1";
defparam ram_block1a5.clk1_input_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "nios_mcu_jtag_uart_0:jtag_uart_0|nios_mcu_jtag_uart_0_scfifo_r:the_nios_mcu_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_jr21:auto_generated|a_dpfifo_l011:dpfifo|altsyncram_nio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 6;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 63;
defparam ram_block1a5.port_a_logical_ram_depth = 64;
defparam ram_block1a5.port_a_logical_ram_width = 8;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 6;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 63;
defparam ram_block1a5.port_b_logical_ram_depth = 64;
defparam ram_block1a5.port_b_logical_ram_width = 8;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk1_core_clock_enable = "ena1";
defparam ram_block1a6.clk1_input_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "nios_mcu_jtag_uart_0:jtag_uart_0|nios_mcu_jtag_uart_0_scfifo_r:the_nios_mcu_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_jr21:auto_generated|a_dpfifo_l011:dpfifo|altsyncram_nio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 6;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 63;
defparam ram_block1a6.port_a_logical_ram_depth = 64;
defparam ram_block1a6.port_a_logical_ram_width = 8;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 6;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 63;
defparam ram_block1a6.port_b_logical_ram_depth = 64;
defparam ram_block1a6.port_b_logical_ram_width = 8;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk1_core_clock_enable = "ena1";
defparam ram_block1a7.clk1_input_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "nios_mcu_jtag_uart_0:jtag_uart_0|nios_mcu_jtag_uart_0_scfifo_r:the_nios_mcu_jtag_uart_0_scfifo_r|scfifo:rfifo|scfifo_jr21:auto_generated|a_dpfifo_l011:dpfifo|altsyncram_nio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 6;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 63;
defparam ram_block1a7.port_a_logical_ram_depth = 64;
defparam ram_block1a7.port_a_logical_ram_width = 8;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 6;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 63;
defparam ram_block1a7.port_b_logical_ram_depth = 64;
defparam ram_block1a7.port_b_logical_ram_width = 8;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

endmodule

module nios_mcu_cntr_1ob (
	r_sync_rst,
	fifo_rd,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	fifo_rd;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5AAF;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout());
defparam counter_comb_bita5.lut_mask = 16'h5A5A;
defparam counter_comb_bita5.sum_lutc_input = "cin";

endmodule

module nios_mcu_cntr_1ob_1 (
	r_sync_rst,
	wr_rfifo,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	wr_rfifo;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5AAF;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout());
defparam counter_comb_bita5.lut_mask = 16'h5A5A;
defparam counter_comb_bita5.sum_lutc_input = "cin";

endmodule

module nios_mcu_nios_mcu_jtag_uart_0_scfifo_w (
	q_b_7,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	d_writedata_0,
	r_sync_rst,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	b_non_empty,
	r_val,
	fifo_wr,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	b_full,
	counter_reg_bit_5,
	counter_reg_bit_4,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_7;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
input 	d_writedata_0;
input 	r_sync_rst;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	d_writedata_6;
input 	d_writedata_7;
output 	b_non_empty;
input 	r_val;
input 	fifo_wr;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	b_full;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nios_mcu_scfifo_2 wfifo(
	.q({q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.data({d_writedata_7,d_writedata_6,d_writedata_5,d_writedata_4,d_writedata_3,d_writedata_2,d_writedata_1,d_writedata_0}),
	.r_sync_rst(r_sync_rst),
	.b_non_empty(b_non_empty),
	.r_val(r_val),
	.wrreq(fifo_wr),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.b_full(b_full),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.clock(clk_clk));

endmodule

module nios_mcu_scfifo_2 (
	q,
	data,
	r_sync_rst,
	b_non_empty,
	r_val,
	wrreq,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	b_full,
	counter_reg_bit_5,
	counter_reg_bit_4,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	[7:0] data;
input 	r_sync_rst;
output 	b_non_empty;
input 	r_val;
input 	wrreq;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	b_full;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nios_mcu_scfifo_jr21_1 auto_generated(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.r_sync_rst(r_sync_rst),
	.b_non_empty(b_non_empty),
	.r_val(r_val),
	.wrreq(wrreq),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.b_full(b_full),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.clock(clock));

endmodule

module nios_mcu_scfifo_jr21_1 (
	q,
	data,
	r_sync_rst,
	b_non_empty,
	r_val,
	wrreq,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	b_full,
	counter_reg_bit_5,
	counter_reg_bit_4,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	[7:0] data;
input 	r_sync_rst;
output 	b_non_empty;
input 	r_val;
input 	wrreq;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	b_full;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nios_mcu_a_dpfifo_l011_1 dpfifo(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.r_sync_rst(r_sync_rst),
	.b_non_empty(b_non_empty),
	.r_val(r_val),
	.wreq(wrreq),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.b_full(b_full),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.clock(clock));

endmodule

module nios_mcu_a_dpfifo_l011_1 (
	q,
	data,
	r_sync_rst,
	b_non_empty,
	r_val,
	wreq,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	b_full,
	counter_reg_bit_5,
	counter_reg_bit_4,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	[7:0] data;
input 	r_sync_rst;
output 	b_non_empty;
input 	r_val;
input 	wreq;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	b_full;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \wr_ptr|counter_reg_bit[5]~q ;
wire \rd_ptr_count|counter_reg_bit[0]~q ;
wire \rd_ptr_count|counter_reg_bit[1]~q ;
wire \rd_ptr_count|counter_reg_bit[2]~q ;
wire \rd_ptr_count|counter_reg_bit[3]~q ;
wire \rd_ptr_count|counter_reg_bit[4]~q ;
wire \rd_ptr_count|counter_reg_bit[5]~q ;


nios_mcu_cntr_1ob_3 wr_ptr(
	.r_sync_rst(r_sync_rst),
	.fifo_wr(wreq),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\wr_ptr|counter_reg_bit[5]~q ),
	.clock(clock));

nios_mcu_cntr_1ob_2 rd_ptr_count(
	.r_sync_rst(r_sync_rst),
	.r_val(r_val),
	.counter_reg_bit_0(\rd_ptr_count|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_count|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_count|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_count|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\rd_ptr_count|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\rd_ptr_count|counter_reg_bit[5]~q ),
	.clock(clock));

nios_mcu_altsyncram_nio1_1 FIFOram(
	.q_b({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data_a({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.clocken1(r_val),
	.wren_a(wreq),
	.address_a({\wr_ptr|counter_reg_bit[5]~q ,\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.address_b({\rd_ptr_count|counter_reg_bit[5]~q ,\rd_ptr_count|counter_reg_bit[4]~q ,\rd_ptr_count|counter_reg_bit[3]~q ,\rd_ptr_count|counter_reg_bit[2]~q ,\rd_ptr_count|counter_reg_bit[1]~q ,\rd_ptr_count|counter_reg_bit[0]~q }),
	.clock0(clock),
	.clock1(clock));

nios_mcu_a_fefifo_7cf_1 fifo_state(
	.r_sync_rst(r_sync_rst),
	.b_non_empty1(b_non_empty),
	.r_val(r_val),
	.wreq(wreq),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.b_full1(b_full),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.clock(clock));

endmodule

module nios_mcu_a_fefifo_7cf_1 (
	r_sync_rst,
	b_non_empty1,
	r_val,
	wreq,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	b_full1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
output 	b_non_empty1;
input 	r_val;
input 	wreq;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	b_full1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \_~0_combout ;
wire \b_non_empty~0_combout ;
wire \b_non_empty~1_combout ;
wire \b_non_empty~2_combout ;
wire \b_full~0_combout ;
wire \b_full~1_combout ;
wire \b_full~2_combout ;


nios_mcu_cntr_do7_1 count_usedw(
	.r_sync_rst(r_sync_rst),
	.updown(wreq),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	._(\_~0_combout ),
	.clock(clock));

cycloneive_lcell_comb \_~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(wreq),
	.datad(r_val),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'h0FF0;
defparam \_~0 .sum_lutc_input = "datac";

dffeas b_non_empty(
	.clk(clock),
	.d(\b_non_empty~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_non_empty1),
	.prn(vcc));
defparam b_non_empty.is_wysiwyg = "true";
defparam b_non_empty.power_up = "low";

dffeas b_full(
	.clk(clock),
	.d(\b_full~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_full1),
	.prn(vcc));
defparam b_full.is_wysiwyg = "true";
defparam b_full.power_up = "low";

cycloneive_lcell_comb \b_non_empty~0 (
	.dataa(counter_reg_bit_2),
	.datab(counter_reg_bit_1),
	.datac(counter_reg_bit_5),
	.datad(counter_reg_bit_4),
	.cin(gnd),
	.combout(\b_non_empty~0_combout ),
	.cout());
defparam \b_non_empty~0 .lut_mask = 16'hFFFE;
defparam \b_non_empty~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_non_empty~1 (
	.dataa(counter_reg_bit_3),
	.datab(\b_non_empty~0_combout ),
	.datac(r_val),
	.datad(counter_reg_bit_0),
	.cin(gnd),
	.combout(\b_non_empty~1_combout ),
	.cout());
defparam \b_non_empty~1 .lut_mask = 16'hEFFF;
defparam \b_non_empty~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_non_empty~2 (
	.dataa(wreq),
	.datab(b_full1),
	.datac(b_non_empty1),
	.datad(\b_non_empty~1_combout ),
	.cin(gnd),
	.combout(\b_non_empty~2_combout ),
	.cout());
defparam \b_non_empty~2 .lut_mask = 16'hFFFE;
defparam \b_non_empty~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_full~0 (
	.dataa(wreq),
	.datab(b_non_empty1),
	.datac(counter_reg_bit_5),
	.datad(counter_reg_bit_4),
	.cin(gnd),
	.combout(\b_full~0_combout ),
	.cout());
defparam \b_full~0 .lut_mask = 16'hFFFE;
defparam \b_full~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_full~1 (
	.dataa(counter_reg_bit_3),
	.datab(counter_reg_bit_0),
	.datac(counter_reg_bit_2),
	.datad(counter_reg_bit_1),
	.cin(gnd),
	.combout(\b_full~1_combout ),
	.cout());
defparam \b_full~1 .lut_mask = 16'hFFFE;
defparam \b_full~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_full~2 (
	.dataa(b_full1),
	.datab(\b_full~0_combout ),
	.datac(\b_full~1_combout ),
	.datad(r_val),
	.cin(gnd),
	.combout(\b_full~2_combout ),
	.cout());
defparam \b_full~2 .lut_mask = 16'hFEFF;
defparam \b_full~2 .sum_lutc_input = "datac";

endmodule

module nios_mcu_cntr_do7_1 (
	r_sync_rst,
	updown,
	counter_reg_bit_3,
	counter_reg_bit_0,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	_,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	updown;
output 	counter_reg_bit_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
input 	_;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita0~combout ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;
wire \counter_comb_bita4~combout ;


dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A6F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5A6F;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout());
defparam counter_comb_bita5.lut_mask = 16'h5A5A;
defparam counter_comb_bita5.sum_lutc_input = "cin";

endmodule

module nios_mcu_altsyncram_nio1_1 (
	q_b,
	data_a,
	clocken1,
	wren_a,
	address_a,
	address_b,
	clock0,
	clock1)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q_b;
input 	[7:0] data_a;
input 	clocken1;
input 	wren_a;
input 	[5:0] address_a;
input 	[5:0] address_b;
input 	clock0;
input 	clock1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk1_core_clock_enable = "ena1";
defparam ram_block1a7.clk1_input_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "nios_mcu_jtag_uart_0:jtag_uart_0|nios_mcu_jtag_uart_0_scfifo_w:the_nios_mcu_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_jr21:auto_generated|a_dpfifo_l011:dpfifo|altsyncram_nio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 6;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 63;
defparam ram_block1a7.port_a_logical_ram_depth = 64;
defparam ram_block1a7.port_a_logical_ram_width = 8;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 6;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 63;
defparam ram_block1a7.port_b_logical_ram_depth = 64;
defparam ram_block1a7.port_b_logical_ram_width = 8;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk1_core_clock_enable = "ena1";
defparam ram_block1a0.clk1_input_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "nios_mcu_jtag_uart_0:jtag_uart_0|nios_mcu_jtag_uart_0_scfifo_w:the_nios_mcu_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_jr21:auto_generated|a_dpfifo_l011:dpfifo|altsyncram_nio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 6;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 63;
defparam ram_block1a0.port_a_logical_ram_depth = 64;
defparam ram_block1a0.port_a_logical_ram_width = 8;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 6;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 63;
defparam ram_block1a0.port_b_logical_ram_depth = 64;
defparam ram_block1a0.port_b_logical_ram_width = 8;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cycloneive_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk1_core_clock_enable = "ena1";
defparam ram_block1a1.clk1_input_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "nios_mcu_jtag_uart_0:jtag_uart_0|nios_mcu_jtag_uart_0_scfifo_w:the_nios_mcu_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_jr21:auto_generated|a_dpfifo_l011:dpfifo|altsyncram_nio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 6;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 63;
defparam ram_block1a1.port_a_logical_ram_depth = 64;
defparam ram_block1a1.port_a_logical_ram_width = 8;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 6;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 63;
defparam ram_block1a1.port_b_logical_ram_depth = 64;
defparam ram_block1a1.port_b_logical_ram_width = 8;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cycloneive_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk1_core_clock_enable = "ena1";
defparam ram_block1a2.clk1_input_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "nios_mcu_jtag_uart_0:jtag_uart_0|nios_mcu_jtag_uart_0_scfifo_w:the_nios_mcu_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_jr21:auto_generated|a_dpfifo_l011:dpfifo|altsyncram_nio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 6;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 63;
defparam ram_block1a2.port_a_logical_ram_depth = 64;
defparam ram_block1a2.port_a_logical_ram_width = 8;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 6;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 63;
defparam ram_block1a2.port_b_logical_ram_depth = 64;
defparam ram_block1a2.port_b_logical_ram_width = 8;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cycloneive_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk1_core_clock_enable = "ena1";
defparam ram_block1a3.clk1_input_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "nios_mcu_jtag_uart_0:jtag_uart_0|nios_mcu_jtag_uart_0_scfifo_w:the_nios_mcu_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_jr21:auto_generated|a_dpfifo_l011:dpfifo|altsyncram_nio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 6;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 63;
defparam ram_block1a3.port_a_logical_ram_depth = 64;
defparam ram_block1a3.port_a_logical_ram_width = 8;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 6;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 63;
defparam ram_block1a3.port_b_logical_ram_depth = 64;
defparam ram_block1a3.port_b_logical_ram_width = 8;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cycloneive_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk1_core_clock_enable = "ena1";
defparam ram_block1a4.clk1_input_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "nios_mcu_jtag_uart_0:jtag_uart_0|nios_mcu_jtag_uart_0_scfifo_w:the_nios_mcu_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_jr21:auto_generated|a_dpfifo_l011:dpfifo|altsyncram_nio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 6;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 63;
defparam ram_block1a4.port_a_logical_ram_depth = 64;
defparam ram_block1a4.port_a_logical_ram_width = 8;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 6;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 63;
defparam ram_block1a4.port_b_logical_ram_depth = 64;
defparam ram_block1a4.port_b_logical_ram_width = 8;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk1_core_clock_enable = "ena1";
defparam ram_block1a5.clk1_input_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "nios_mcu_jtag_uart_0:jtag_uart_0|nios_mcu_jtag_uart_0_scfifo_w:the_nios_mcu_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_jr21:auto_generated|a_dpfifo_l011:dpfifo|altsyncram_nio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 6;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 63;
defparam ram_block1a5.port_a_logical_ram_depth = 64;
defparam ram_block1a5.port_a_logical_ram_width = 8;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 6;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 63;
defparam ram_block1a5.port_b_logical_ram_depth = 64;
defparam ram_block1a5.port_b_logical_ram_width = 8;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk1_core_clock_enable = "ena1";
defparam ram_block1a6.clk1_input_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "nios_mcu_jtag_uart_0:jtag_uart_0|nios_mcu_jtag_uart_0_scfifo_w:the_nios_mcu_jtag_uart_0_scfifo_w|scfifo:wfifo|scfifo_jr21:auto_generated|a_dpfifo_l011:dpfifo|altsyncram_nio1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 6;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 63;
defparam ram_block1a6.port_a_logical_ram_depth = 64;
defparam ram_block1a6.port_a_logical_ram_width = 8;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 6;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 63;
defparam ram_block1a6.port_b_logical_ram_depth = 64;
defparam ram_block1a6.port_b_logical_ram_width = 8;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

endmodule

module nios_mcu_cntr_1ob_2 (
	r_sync_rst,
	r_val,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	r_val;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5AAF;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout());
defparam counter_comb_bita5.lut_mask = 16'h5A5A;
defparam counter_comb_bita5.sum_lutc_input = "cin";

endmodule

module nios_mcu_cntr_1ob_3 (
	r_sync_rst,
	fifo_wr,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	fifo_wr;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout(\counter_comb_bita4~COUT ));
defparam counter_comb_bita4.lut_mask = 16'h5AAF;
defparam counter_comb_bita4.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita5(
	.dataa(counter_reg_bit_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.combout(\counter_comb_bita5~combout ),
	.cout());
defparam counter_comb_bita5.lut_mask = 16'h5A5A;
defparam counter_comb_bita5.sum_lutc_input = "cin";

endmodule

module nios_mcu_nios_mcu_mm_interconnect_0 (
	W_alu_result_12,
	W_alu_result_15,
	W_alu_result_14,
	W_alu_result_13,
	W_alu_result_11,
	W_alu_result_10,
	W_alu_result_9,
	W_alu_result_8,
	W_alu_result_7,
	W_alu_result_6,
	W_alu_result_5,
	W_alu_result_4,
	W_alu_result_3,
	W_alu_result_2,
	q_b_22,
	q_b_23,
	q_a_11,
	q_b_11,
	q_a_13,
	q_b_13,
	q_a_16,
	q_b_16,
	q_b_12,
	q_a_1,
	q_a_3,
	q_a_5,
	q_a_4,
	q_b_14,
	q_a_15,
	q_b_15,
	q_b_18,
	q_b_17,
	q_b_10,
	q_b_9,
	q_b_8,
	q_a_21,
	q_b_21,
	q_a_19,
	q_b_19,
	q_a_20,
	q_b_20,
	readdata_0,
	d_writedata_24,
	d_writedata_25,
	d_writedata_26,
	readdata_1,
	readdata_3,
	readdata_2,
	d_writedata_27,
	d_writedata_28,
	d_writedata_29,
	d_writedata_30,
	d_writedata_31,
	d_writedata_0,
	r_sync_rst,
	Equal1,
	rst1,
	mem_used_1,
	always0,
	d_write,
	write_accepted,
	wait_latency_counter_1,
	wait_latency_counter_0,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	read_latency_shift_reg_0,
	d_read,
	read_latency_shift_reg,
	m0_write,
	mem_73_0,
	mem_55_0,
	read_latency_shift_reg_01,
	read_latency_shift_reg_02,
	WideOr1,
	read_latency_shift_reg_03,
	read_latency_shift_reg_04,
	WideOr11,
	Equal3,
	src_channel_4,
	mem_used_11,
	saved_grant_0,
	waitrequest,
	mem_used_12,
	av_waitrequest,
	mem_used_13,
	Equal2,
	dRead,
	always2,
	m0_read,
	m0_read1,
	sReadCountPipelined_0,
	nios_cpu_data_master_waitrequest,
	F_pc_10,
	F_pc_9,
	F_pc_8,
	F_pc_7,
	F_pc_6,
	F_pc_5,
	F_pc_4,
	F_pc_3,
	F_pc_2,
	F_pc_1,
	F_pc_0,
	F_pc_13,
	F_pc_12,
	F_pc_11,
	i_read,
	WideOr12,
	Equal21,
	rf_source_valid,
	hbreak_enabled,
	WideOr13,
	av_readdata_pre_0,
	av_readdata_pre_01,
	av_readdata_pre_02,
	src0_valid,
	av_readdata_pre_03,
	av_readdata_pre_22,
	read_latency_shift_reg_05,
	src1_valid,
	av_readdata_pre_23,
	av_readdata_pre_24,
	av_readdata_pre_25,
	av_readdata_pre_26,
	src_payload,
	av_readdata_pre_11,
	src_payload1,
	av_readdata_pre_13,
	src_payload2,
	av_readdata_pre_16,
	av_readdata_pre_12,
	src_payload3,
	av_readdata_pre_1,
	src_payload4,
	av_readdata_pre_3,
	av_readdata_pre_2,
	src_payload5,
	av_readdata_pre_5,
	src_payload6,
	av_readdata_pre_4,
	av_readdata_pre_14,
	src_payload7,
	av_readdata_pre_15,
	av_readdata_pre_18,
	av_readdata_pre_17,
	av_readdata_pre_10,
	av_readdata_pre_9,
	av_readdata_pre_8,
	av_readdata_pre_7,
	av_readdata_pre_6,
	src_payload8,
	av_readdata_pre_21,
	src_payload9,
	av_readdata_pre_19,
	src_payload10,
	av_readdata_pre_20,
	src_data_46,
	av_readdata_pre_110,
	av_readdata_pre_111,
	av_readdata_pre_112,
	av_readdata_pre_27,
	av_readdata_pre_28,
	av_readdata_pre_29,
	av_readdata_pre_31,
	av_readdata_pre_32,
	av_readdata_pre_33,
	av_readdata_pre_41,
	av_readdata_pre_42,
	av_readdata_pre_43,
	av_readdata_pre_51,
	av_readdata_pre_52,
	av_readdata_pre_53,
	av_readdata_pre_61,
	av_readdata_pre_62,
	av_readdata_pre_63,
	av_readdata_pre_71,
	av_readdata_pre_72,
	av_readdata_pre_73,
	b_full,
	src_data_8,
	ReadData_0,
	read_0,
	av_readdata_0,
	d_byteenable_0,
	readdata_01,
	av_readdata_9,
	av_readdata_8,
	readdata_22,
	d_writedata_22,
	d_byteenable_2,
	readdata_23,
	d_writedata_23,
	readdata_24,
	d_byteenable_3,
	readdata_25,
	readdata_26,
	d_writedata_11,
	d_byteenable_1,
	readdata_11,
	d_writedata_13,
	readdata_13,
	d_writedata_16,
	readdata_16,
	readdata_12,
	d_writedata_12,
	readdata_5,
	readdata_4,
	d_writedata_14,
	readdata_14,
	d_writedata_15,
	readdata_15,
	d_writedata_18,
	readdata_18,
	src_data_12,
	av_readdata_pre_271,
	av_readdata_pre_281,
	av_readdata_pre_291,
	av_readdata_pre_30,
	av_readdata_pre_311,
	d_writedata_17,
	readdata_17,
	src_data_11,
	src_data_10,
	src_data_9,
	readdata_10,
	d_writedata_10,
	readdata_9,
	d_writedata_9,
	readdata_8,
	d_writedata_8,
	readdata_7,
	readdata_6,
	d_writedata_21,
	readdata_21,
	src_data_15,
	d_writedata_19,
	readdata_19,
	d_writedata_20,
	readdata_20,
	src_data_14,
	src_data_13,
	ReadData_1,
	av_readdata_1,
	readdata_110,
	ReadData_2,
	av_readdata_2,
	readdata_27,
	ReadData_3,
	av_readdata_3,
	readdata_31,
	ReadData_4,
	av_readdata_4,
	readdata_41,
	ReadData_5,
	av_readdata_5,
	readdata_51,
	ReadData_6,
	av_readdata_6,
	readdata_61,
	ReadData_7,
	av_readdata_7,
	readdata_71,
	b_non_empty,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	src_payload11,
	src_payload12,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_32,
	ReadData_8,
	src_data_16,
	counter_reg_bit_31,
	counter_reg_bit_01,
	counter_reg_bit_21,
	counter_reg_bit_11,
	b_full1,
	counter_reg_bit_51,
	counter_reg_bit_41,
	ReadData_12,
	src_data_20,
	readdata_271,
	readdata_28,
	readdata_29,
	readdata_30,
	readdata_311,
	ReadData_11,
	src_data_19,
	ReadData_10,
	ac,
	src_data_18,
	ReadData_9,
	src_data_17,
	ReadData_15,
	rvalid,
	src_data_23,
	ReadData_14,
	woverflow,
	src_data_22,
	ReadData_13,
	src_data_21,
	src_payload13,
	ReadData_16,
	av_readdata_pre_241,
	av_readdata_pre_312,
	av_readdata_pre_301,
	av_readdata_pre_292,
	av_readdata_pre_282,
	av_readdata_pre_272,
	av_readdata_pre_261,
	av_readdata_pre_251,
	src_payload14,
	ReadData_20,
	ReadData_19,
	ReadData_18,
	ReadData_17,
	ReadData_23,
	ReadData_22,
	ReadData_21,
	src_payload15,
	ReadData_24,
	ReadData_31,
	ReadData_30,
	ReadData_29,
	ReadData_28,
	ReadData_27,
	ReadData_26,
	ReadData_25,
	src_payload16,
	src_data_34,
	src_payload17,
	src_payload18,
	src_data_35,
	src_payload19,
	src_payload20,
	src_payload21,
	src_data_33,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32,
	src_payload33,
	src_payload34,
	src_payload35,
	src_payload36,
	src_payload37,
	src_payload38,
	src_payload39,
	src_payload40,
	src_payload41,
	src_payload42,
	src_payload43,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_12;
input 	W_alu_result_15;
input 	W_alu_result_14;
input 	W_alu_result_13;
input 	W_alu_result_11;
input 	W_alu_result_10;
input 	W_alu_result_9;
input 	W_alu_result_8;
input 	W_alu_result_7;
input 	W_alu_result_6;
input 	W_alu_result_5;
input 	W_alu_result_4;
input 	W_alu_result_3;
input 	W_alu_result_2;
input 	q_b_22;
input 	q_b_23;
input 	q_a_11;
input 	q_b_11;
input 	q_a_13;
input 	q_b_13;
input 	q_a_16;
input 	q_b_16;
input 	q_b_12;
input 	q_a_1;
input 	q_a_3;
input 	q_a_5;
input 	q_a_4;
input 	q_b_14;
input 	q_a_15;
input 	q_b_15;
input 	q_b_18;
input 	q_b_17;
input 	q_b_10;
input 	q_b_9;
input 	q_b_8;
input 	q_a_21;
input 	q_b_21;
input 	q_a_19;
input 	q_b_19;
input 	q_a_20;
input 	q_b_20;
input 	readdata_0;
input 	d_writedata_24;
input 	d_writedata_25;
input 	d_writedata_26;
input 	readdata_1;
input 	readdata_3;
input 	readdata_2;
input 	d_writedata_27;
input 	d_writedata_28;
input 	d_writedata_29;
input 	d_writedata_30;
input 	d_writedata_31;
input 	d_writedata_0;
input 	r_sync_rst;
output 	Equal1;
input 	rst1;
output 	mem_used_1;
input 	always0;
input 	d_write;
output 	write_accepted;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	d_writedata_6;
input 	d_writedata_7;
output 	read_latency_shift_reg_0;
input 	d_read;
output 	read_latency_shift_reg;
output 	m0_write;
output 	mem_73_0;
output 	mem_55_0;
output 	read_latency_shift_reg_01;
output 	read_latency_shift_reg_02;
output 	WideOr1;
output 	read_latency_shift_reg_03;
output 	read_latency_shift_reg_04;
output 	WideOr11;
output 	Equal3;
output 	src_channel_4;
output 	mem_used_11;
output 	saved_grant_0;
input 	waitrequest;
output 	mem_used_12;
input 	av_waitrequest;
output 	mem_used_13;
output 	Equal2;
input 	dRead;
output 	always2;
output 	m0_read;
output 	m0_read1;
input 	sReadCountPipelined_0;
output 	nios_cpu_data_master_waitrequest;
input 	F_pc_10;
input 	F_pc_9;
input 	F_pc_8;
input 	F_pc_7;
input 	F_pc_6;
input 	F_pc_5;
input 	F_pc_4;
input 	F_pc_3;
input 	F_pc_2;
input 	F_pc_1;
input 	F_pc_0;
input 	F_pc_13;
input 	F_pc_12;
input 	F_pc_11;
input 	i_read;
output 	WideOr12;
input 	Equal21;
output 	rf_source_valid;
input 	hbreak_enabled;
output 	WideOr13;
output 	av_readdata_pre_0;
output 	av_readdata_pre_01;
output 	av_readdata_pre_02;
output 	src0_valid;
output 	av_readdata_pre_03;
output 	av_readdata_pre_22;
output 	read_latency_shift_reg_05;
output 	src1_valid;
output 	av_readdata_pre_23;
output 	av_readdata_pre_24;
output 	av_readdata_pre_25;
output 	av_readdata_pre_26;
output 	src_payload;
output 	av_readdata_pre_11;
output 	src_payload1;
output 	av_readdata_pre_13;
output 	src_payload2;
output 	av_readdata_pre_16;
output 	av_readdata_pre_12;
output 	src_payload3;
output 	av_readdata_pre_1;
output 	src_payload4;
output 	av_readdata_pre_3;
output 	av_readdata_pre_2;
output 	src_payload5;
output 	av_readdata_pre_5;
output 	src_payload6;
output 	av_readdata_pre_4;
output 	av_readdata_pre_14;
output 	src_payload7;
output 	av_readdata_pre_15;
output 	av_readdata_pre_18;
output 	av_readdata_pre_17;
output 	av_readdata_pre_10;
output 	av_readdata_pre_9;
output 	av_readdata_pre_8;
output 	av_readdata_pre_7;
output 	av_readdata_pre_6;
output 	src_payload8;
output 	av_readdata_pre_21;
output 	src_payload9;
output 	av_readdata_pre_19;
output 	src_payload10;
output 	av_readdata_pre_20;
output 	src_data_46;
output 	av_readdata_pre_110;
output 	av_readdata_pre_111;
output 	av_readdata_pre_112;
output 	av_readdata_pre_27;
output 	av_readdata_pre_28;
output 	av_readdata_pre_29;
output 	av_readdata_pre_31;
output 	av_readdata_pre_32;
output 	av_readdata_pre_33;
output 	av_readdata_pre_41;
output 	av_readdata_pre_42;
output 	av_readdata_pre_43;
output 	av_readdata_pre_51;
output 	av_readdata_pre_52;
output 	av_readdata_pre_53;
output 	av_readdata_pre_61;
output 	av_readdata_pre_62;
output 	av_readdata_pre_63;
output 	av_readdata_pre_71;
output 	av_readdata_pre_72;
output 	av_readdata_pre_73;
input 	b_full;
output 	src_data_8;
input 	ReadData_0;
input 	read_0;
input 	av_readdata_0;
input 	d_byteenable_0;
input 	readdata_01;
input 	av_readdata_9;
input 	av_readdata_8;
input 	readdata_22;
input 	d_writedata_22;
input 	d_byteenable_2;
input 	readdata_23;
input 	d_writedata_23;
input 	readdata_24;
input 	d_byteenable_3;
input 	readdata_25;
input 	readdata_26;
input 	d_writedata_11;
input 	d_byteenable_1;
input 	readdata_11;
input 	d_writedata_13;
input 	readdata_13;
input 	d_writedata_16;
input 	readdata_16;
input 	readdata_12;
input 	d_writedata_12;
input 	readdata_5;
input 	readdata_4;
input 	d_writedata_14;
input 	readdata_14;
input 	d_writedata_15;
input 	readdata_15;
input 	d_writedata_18;
input 	readdata_18;
output 	src_data_12;
output 	av_readdata_pre_271;
output 	av_readdata_pre_281;
output 	av_readdata_pre_291;
output 	av_readdata_pre_30;
output 	av_readdata_pre_311;
input 	d_writedata_17;
input 	readdata_17;
output 	src_data_11;
output 	src_data_10;
output 	src_data_9;
input 	readdata_10;
input 	d_writedata_10;
input 	readdata_9;
input 	d_writedata_9;
input 	readdata_8;
input 	d_writedata_8;
input 	readdata_7;
input 	readdata_6;
input 	d_writedata_21;
input 	readdata_21;
output 	src_data_15;
input 	d_writedata_19;
input 	readdata_19;
input 	d_writedata_20;
input 	readdata_20;
output 	src_data_14;
output 	src_data_13;
input 	ReadData_1;
input 	av_readdata_1;
input 	readdata_110;
input 	ReadData_2;
input 	av_readdata_2;
input 	readdata_27;
input 	ReadData_3;
input 	av_readdata_3;
input 	readdata_31;
input 	ReadData_4;
input 	av_readdata_4;
input 	readdata_41;
input 	ReadData_5;
input 	av_readdata_5;
input 	readdata_51;
input 	ReadData_6;
input 	av_readdata_6;
input 	readdata_61;
input 	ReadData_7;
input 	av_readdata_7;
input 	readdata_71;
input 	b_non_empty;
input 	counter_reg_bit_5;
input 	counter_reg_bit_4;
input 	counter_reg_bit_3;
input 	counter_reg_bit_2;
input 	counter_reg_bit_1;
input 	counter_reg_bit_0;
output 	src_payload11;
output 	src_payload12;
output 	src_data_38;
output 	src_data_39;
output 	src_data_40;
output 	src_data_41;
output 	src_data_42;
output 	src_data_43;
output 	src_data_44;
output 	src_data_45;
output 	src_data_32;
input 	ReadData_8;
output 	src_data_16;
input 	counter_reg_bit_31;
input 	counter_reg_bit_01;
input 	counter_reg_bit_21;
input 	counter_reg_bit_11;
input 	b_full1;
input 	counter_reg_bit_51;
input 	counter_reg_bit_41;
input 	ReadData_12;
output 	src_data_20;
input 	readdata_271;
input 	readdata_28;
input 	readdata_29;
input 	readdata_30;
input 	readdata_311;
input 	ReadData_11;
output 	src_data_19;
input 	ReadData_10;
input 	ac;
output 	src_data_18;
input 	ReadData_9;
output 	src_data_17;
input 	ReadData_15;
input 	rvalid;
output 	src_data_23;
input 	ReadData_14;
input 	woverflow;
output 	src_data_22;
input 	ReadData_13;
output 	src_data_21;
output 	src_payload13;
input 	ReadData_16;
output 	av_readdata_pre_241;
output 	av_readdata_pre_312;
output 	av_readdata_pre_301;
output 	av_readdata_pre_292;
output 	av_readdata_pre_282;
output 	av_readdata_pre_272;
output 	av_readdata_pre_261;
output 	av_readdata_pre_251;
output 	src_payload14;
input 	ReadData_20;
input 	ReadData_19;
input 	ReadData_18;
input 	ReadData_17;
input 	ReadData_23;
input 	ReadData_22;
input 	ReadData_21;
output 	src_payload15;
input 	ReadData_24;
input 	ReadData_31;
input 	ReadData_30;
input 	ReadData_29;
input 	ReadData_28;
input 	ReadData_27;
input 	ReadData_26;
input 	ReadData_25;
output 	src_payload16;
output 	src_data_34;
output 	src_payload17;
output 	src_payload18;
output 	src_data_35;
output 	src_payload19;
output 	src_payload20;
output 	src_payload21;
output 	src_data_33;
output 	src_payload22;
output 	src_payload23;
output 	src_payload24;
output 	src_payload25;
output 	src_payload26;
output 	src_payload27;
output 	src_payload28;
output 	src_payload29;
output 	src_payload30;
output 	src_payload31;
output 	src_payload32;
output 	src_payload33;
output 	src_payload34;
output 	src_payload35;
output 	src_payload36;
output 	src_payload37;
output 	src_payload38;
output 	src_payload39;
output 	src_payload40;
output 	src_payload41;
output 	src_payload42;
output 	src_payload43;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[16]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[20]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[19]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[18]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[17]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[22]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[21]~q ;
wire \nios_cpu_data_master_translator|read_accepted~q ;
wire \router|Equal1~4_combout ;
wire \pio_0_s1_translator|wait_latency_counter[1]~0_combout ;
wire \router|Equal0~0_combout ;
wire \cmd_demux|sink_ready~0_combout ;
wire \nios_cpu_debug_mem_slave_agent_rsp_fifo|write~0_combout ;
wire \cmd_demux|WideOr0~0_combout ;
wire \pio_0_s1_translator|read_latency_shift_reg~0_combout ;
wire \nios_cpu_data_master_translator|uav_read~0_combout ;
wire \avalonslave_0_avalon_slave_0_1_agent_rsp_fifo|mem_used[1]~q ;
wire \cmd_demux|sink_ready~2_combout ;
wire \cmd_demux|WideOr0~1_combout ;
wire \pio_0_s1_translator|read_latency_shift_reg~1_combout ;
wire \cmd_mux_002|saved_grant[1]~q ;
wire \nios_cpu_debug_mem_slave_agent|rf_source_valid~0_combout ;
wire \nios_cpu_instruction_master_translator|read_accepted~q ;
wire \nios_cpu_debug_mem_slave_agent_rsp_fifo|mem~1_combout ;
wire \onchip_ram_s1_translator|read_latency_shift_reg~0_combout ;
wire \router_001|Equal0~0_combout ;
wire \cmd_demux_001|src0_valid~0_combout ;
wire \cmd_demux|src2_valid~0_combout ;
wire \jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg~1_combout ;
wire \avalonslave_0_avalon_slave_0_1_translator|read_latency_shift_reg~0_combout ;
wire \onchip_ram_s2_translator|read_latency_shift_reg~0_combout ;
wire \router_001|Equal0~1_combout ;
wire \onchip_ram_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[8]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[8]~q ;
wire \onchip_ram_s1_translator|read_latency_shift_reg~1_combout ;
wire \avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[12]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[12]~q ;
wire \avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[11]~q ;
wire \avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[10]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[10]~q ;
wire \avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[9]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[9]~q ;
wire \avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[15]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[15]~q ;
wire \avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[14]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[14]~q ;
wire \avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[13]~q ;
wire \jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[13]~q ;
wire \avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[16]~q ;
wire \avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[20]~q ;
wire \avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[19]~q ;
wire \avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[18]~q ;
wire \avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[17]~q ;
wire \avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[23]~q ;
wire \avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[22]~q ;
wire \avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[21]~q ;


nios_mcu_altera_avalon_sc_fifo_4 onchip_ram_s2_agent_rsp_fifo(
	.reset(r_sync_rst),
	.read_latency_shift_reg(read_latency_shift_reg),
	.read_latency_shift_reg_0(read_latency_shift_reg_04),
	.src_channel_4(src_channel_4),
	.mem_used_1(mem_used_11),
	.read_latency_shift_reg1(\onchip_ram_s2_translator|read_latency_shift_reg~0_combout ),
	.clk(clk_clk));

nios_mcu_altera_avalon_sc_fifo_5 pio_0_s1_agent_rsp_fifo(
	.W_alu_result_4(W_alu_result_4),
	.reset(r_sync_rst),
	.Equal1(Equal1),
	.mem_used_1(mem_used_1),
	.read_latency_shift_reg_0(read_latency_shift_reg_0),
	.read_latency_shift_reg(read_latency_shift_reg),
	.wait_latency_counter_1(\pio_0_s1_translator|wait_latency_counter[1]~0_combout ),
	.read_latency_shift_reg1(\pio_0_s1_translator|read_latency_shift_reg~1_combout ),
	.clk(clk_clk));

nios_mcu_altera_merlin_slave_agent_5 pio_0_s1_agent(
	.d_write(d_write),
	.write_accepted(write_accepted),
	.m0_write(m0_write));

nios_mcu_altera_avalon_sc_fifo_2 nios_cpu_debug_mem_slave_agent_rsp_fifo(
	.reset(r_sync_rst),
	.mem_73_0(mem_73_0),
	.mem_55_0(mem_55_0),
	.read_latency_shift_reg_0(read_latency_shift_reg_01),
	.waitrequest(waitrequest),
	.mem_used_1(mem_used_12),
	.write(\nios_cpu_debug_mem_slave_agent_rsp_fifo|write~0_combout ),
	.saved_grant_1(\cmd_mux_002|saved_grant[1]~q ),
	.rf_source_valid(\nios_cpu_debug_mem_slave_agent|rf_source_valid~0_combout ),
	.read_accepted(\nios_cpu_instruction_master_translator|read_accepted~q ),
	.i_read(i_read),
	.mem(\nios_cpu_debug_mem_slave_agent_rsp_fifo|mem~1_combout ),
	.WideOr1(WideOr12),
	.rf_source_valid1(rf_source_valid),
	.clk(clk_clk));

nios_mcu_altera_merlin_slave_agent_2 nios_cpu_debug_mem_slave_agent(
	.d_read(d_read),
	.read_accepted(\nios_cpu_data_master_translator|read_accepted~q ),
	.saved_grant_0(saved_grant_0),
	.rf_source_valid(\nios_cpu_debug_mem_slave_agent|rf_source_valid~0_combout ),
	.mem(\nios_cpu_debug_mem_slave_agent_rsp_fifo|mem~1_combout ),
	.WideOr1(WideOr12),
	.rf_source_valid1(rf_source_valid));

nios_mcu_altera_avalon_sc_fifo avalonslave_0_avalon_slave_0_1_agent_rsp_fifo(
	.reset(r_sync_rst),
	.rst1(rst1),
	.read_latency_shift_reg_0(read_latency_shift_reg_03),
	.Equal2(Equal2),
	.uav_read(\nios_cpu_data_master_translator|uav_read~0_combout ),
	.mem_used_1(\avalonslave_0_avalon_slave_0_1_agent_rsp_fifo|mem_used[1]~q ),
	.Equal21(Equal21),
	.read_latency_shift_reg(\avalonslave_0_avalon_slave_0_1_translator|read_latency_shift_reg~0_combout ),
	.clk(clk_clk));

nios_mcu_nios_mcu_mm_interconnect_0_cmd_mux_002 cmd_mux_002(
	.W_alu_result_10(W_alu_result_10),
	.W_alu_result_9(W_alu_result_9),
	.W_alu_result_8(W_alu_result_8),
	.W_alu_result_7(W_alu_result_7),
	.W_alu_result_6(W_alu_result_6),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_3(W_alu_result_3),
	.W_alu_result_2(W_alu_result_2),
	.d_writedata_24(d_writedata_24),
	.d_writedata_25(d_writedata_25),
	.d_writedata_26(d_writedata_26),
	.d_writedata_27(d_writedata_27),
	.d_writedata_28(d_writedata_28),
	.d_writedata_29(d_writedata_29),
	.d_writedata_30(d_writedata_30),
	.d_writedata_31(d_writedata_31),
	.d_writedata_0(d_writedata_0),
	.r_sync_rst(r_sync_rst),
	.d_writedata_1(d_writedata_1),
	.d_writedata_2(d_writedata_2),
	.d_writedata_3(d_writedata_3),
	.d_writedata_4(d_writedata_4),
	.d_writedata_5(d_writedata_5),
	.d_writedata_6(d_writedata_6),
	.d_writedata_7(d_writedata_7),
	.saved_grant_0(saved_grant_0),
	.waitrequest(waitrequest),
	.mem_used_1(mem_used_12),
	.F_pc_8(F_pc_8),
	.F_pc_7(F_pc_7),
	.F_pc_6(F_pc_6),
	.F_pc_5(F_pc_5),
	.F_pc_4(F_pc_4),
	.F_pc_3(F_pc_3),
	.F_pc_2(F_pc_2),
	.F_pc_1(F_pc_1),
	.F_pc_0(F_pc_0),
	.saved_grant_1(\cmd_mux_002|saved_grant[1]~q ),
	.src0_valid(\cmd_demux_001|src0_valid~0_combout ),
	.src2_valid(\cmd_demux|src2_valid~0_combout ),
	.WideOr11(WideOr12),
	.hbreak_enabled(hbreak_enabled),
	.src_data_46(src_data_46),
	.d_byteenable_0(d_byteenable_0),
	.d_writedata_22(d_writedata_22),
	.d_byteenable_2(d_byteenable_2),
	.d_writedata_23(d_writedata_23),
	.d_byteenable_3(d_byteenable_3),
	.d_writedata_11(d_writedata_11),
	.d_byteenable_1(d_byteenable_1),
	.d_writedata_13(d_writedata_13),
	.d_writedata_16(d_writedata_16),
	.d_writedata_12(d_writedata_12),
	.d_writedata_14(d_writedata_14),
	.d_writedata_15(d_writedata_15),
	.d_writedata_18(d_writedata_18),
	.d_writedata_17(d_writedata_17),
	.d_writedata_10(d_writedata_10),
	.d_writedata_9(d_writedata_9),
	.d_writedata_8(d_writedata_8),
	.d_writedata_21(d_writedata_21),
	.d_writedata_19(d_writedata_19),
	.d_writedata_20(d_writedata_20),
	.src_payload(src_payload11),
	.src_payload1(src_payload12),
	.src_data_38(src_data_38),
	.src_data_39(src_data_39),
	.src_data_40(src_data_40),
	.src_data_41(src_data_41),
	.src_data_42(src_data_42),
	.src_data_43(src_data_43),
	.src_data_44(src_data_44),
	.src_data_45(src_data_45),
	.src_data_32(src_data_32),
	.src_payload2(src_payload13),
	.src_payload3(src_payload14),
	.src_payload4(src_payload15),
	.src_payload5(src_payload16),
	.src_data_34(src_data_34),
	.src_payload6(src_payload17),
	.src_payload7(src_payload18),
	.src_data_35(src_data_35),
	.src_payload8(src_payload19),
	.src_payload9(src_payload20),
	.src_payload10(src_payload21),
	.src_data_33(src_data_33),
	.src_payload11(src_payload22),
	.src_payload12(src_payload23),
	.src_payload13(src_payload24),
	.src_payload14(src_payload25),
	.src_payload15(src_payload26),
	.src_payload16(src_payload27),
	.src_payload17(src_payload28),
	.src_payload18(src_payload29),
	.src_payload19(src_payload30),
	.src_payload20(src_payload31),
	.src_payload21(src_payload32),
	.src_payload22(src_payload33),
	.src_payload23(src_payload34),
	.src_payload24(src_payload35),
	.src_payload25(src_payload36),
	.src_payload26(src_payload37),
	.src_payload27(src_payload38),
	.src_payload28(src_payload39),
	.src_payload29(src_payload40),
	.src_payload30(src_payload41),
	.src_payload31(src_payload42),
	.src_payload32(src_payload43),
	.clk_clk(clk_clk));

nios_mcu_nios_mcu_mm_interconnect_0_cmd_demux_001 cmd_demux_001(
	.F_pc_9(F_pc_9),
	.read_latency_shift_reg(\onchip_ram_s1_translator|read_latency_shift_reg~0_combout ),
	.Equal0(\router_001|Equal0~0_combout ),
	.src0_valid(\cmd_demux_001|src0_valid~0_combout ));

nios_mcu_nios_mcu_mm_interconnect_0_cmd_demux cmd_demux(
	.W_alu_result_11(W_alu_result_11),
	.rst1(rst1),
	.Equal0(\router|Equal0~0_combout ),
	.Equal3(Equal3),
	.src_channel_4(src_channel_4),
	.mem_used_1(mem_used_11),
	.sink_ready(\cmd_demux|sink_ready~0_combout ),
	.saved_grant_0(saved_grant_0),
	.write(\nios_cpu_debug_mem_slave_agent_rsp_fifo|write~0_combout ),
	.av_waitrequest(av_waitrequest),
	.mem_used_11(mem_used_13),
	.WideOr0(\cmd_demux|WideOr0~0_combout ),
	.Equal2(Equal2),
	.dRead(dRead),
	.always2(always2),
	.mem_used_12(\avalonslave_0_avalon_slave_0_1_agent_rsp_fifo|mem_used[1]~q ),
	.sReadCountPipelined_0(sReadCountPipelined_0),
	.sink_ready1(\cmd_demux|sink_ready~2_combout ),
	.WideOr01(\cmd_demux|WideOr0~1_combout ),
	.src2_valid(\cmd_demux|src2_valid~0_combout ));

nios_mcu_nios_mcu_mm_interconnect_0_router_001 router_001(
	.F_pc_10(F_pc_10),
	.F_pc_9(F_pc_9),
	.F_pc_13(F_pc_13),
	.F_pc_12(F_pc_12),
	.F_pc_11(F_pc_11),
	.Equal0(\router_001|Equal0~0_combout ),
	.Equal01(\router_001|Equal0~1_combout ));

nios_mcu_nios_mcu_mm_interconnect_0_router router(
	.W_alu_result_12(W_alu_result_12),
	.W_alu_result_15(W_alu_result_15),
	.W_alu_result_14(W_alu_result_14),
	.W_alu_result_13(W_alu_result_13),
	.W_alu_result_11(W_alu_result_11),
	.W_alu_result_10(W_alu_result_10),
	.W_alu_result_9(W_alu_result_9),
	.W_alu_result_8(W_alu_result_8),
	.W_alu_result_7(W_alu_result_7),
	.W_alu_result_6(W_alu_result_6),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_3(W_alu_result_3),
	.Equal1(Equal1),
	.Equal11(\router|Equal1~4_combout ),
	.Equal0(\router|Equal0~0_combout ),
	.Equal3(Equal3),
	.src_channel_4(src_channel_4),
	.Equal2(Equal2));

nios_mcu_altera_avalon_sc_fifo_3 onchip_ram_s1_agent_rsp_fifo(
	.reset(r_sync_rst),
	.read_latency_shift_reg(\onchip_ram_s1_translator|read_latency_shift_reg~0_combout ),
	.read_latency_shift_reg_0(read_latency_shift_reg_05),
	.Equal0(\router_001|Equal0~1_combout ),
	.mem_used_1(\onchip_ram_s1_agent_rsp_fifo|mem_used[1]~q ),
	.read_latency_shift_reg1(\onchip_ram_s1_translator|read_latency_shift_reg~1_combout ),
	.clk(clk_clk));

nios_mcu_nios_mcu_mm_interconnect_0_rsp_mux_001 rsp_mux_001(
	.q_a_11(q_a_11),
	.q_a_13(q_a_13),
	.q_a_16(q_a_16),
	.q_a_1(q_a_1),
	.q_a_3(q_a_3),
	.q_a_5(q_a_5),
	.q_a_4(q_a_4),
	.q_a_15(q_a_15),
	.q_a_21(q_a_21),
	.q_a_19(q_a_19),
	.q_a_20(q_a_20),
	.read_latency_shift_reg_0(read_latency_shift_reg_05),
	.src_payload(src_payload),
	.src_payload1(src_payload1),
	.src_payload2(src_payload2),
	.src_payload3(src_payload3),
	.src_payload4(src_payload4),
	.src_payload5(src_payload5),
	.src_payload6(src_payload6),
	.src_payload7(src_payload7),
	.src_payload8(src_payload8),
	.src_payload9(src_payload9),
	.src_payload10(src_payload10));

nios_mcu_nios_mcu_mm_interconnect_0_rsp_mux rsp_mux(
	.q_b_22(q_b_22),
	.q_b_23(q_b_23),
	.q_b_11(q_b_11),
	.q_b_13(q_b_13),
	.q_b_16(q_b_16),
	.q_b_12(q_b_12),
	.q_b_14(q_b_14),
	.q_b_15(q_b_15),
	.q_b_18(q_b_18),
	.q_b_17(q_b_17),
	.q_b_10(q_b_10),
	.q_b_9(q_b_9),
	.q_b_8(q_b_8),
	.q_b_21(q_b_21),
	.q_b_19(q_b_19),
	.q_b_20(q_b_20),
	.av_readdata_pre_16(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[16]~q ),
	.av_readdata_pre_20(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[20]~q ),
	.av_readdata_pre_19(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[19]~q ),
	.av_readdata_pre_18(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[18]~q ),
	.av_readdata_pre_17(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[17]~q ),
	.av_readdata_pre_22(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[22]~q ),
	.av_readdata_pre_21(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[21]~q ),
	.read_latency_shift_reg_0(read_latency_shift_reg_0),
	.mem_73_0(mem_73_0),
	.mem_55_0(mem_55_0),
	.read_latency_shift_reg_01(read_latency_shift_reg_01),
	.read_latency_shift_reg_02(read_latency_shift_reg_02),
	.WideOr11(WideOr1),
	.read_latency_shift_reg_03(read_latency_shift_reg_03),
	.read_latency_shift_reg_04(read_latency_shift_reg_04),
	.WideOr12(WideOr11),
	.WideOr13(WideOr13),
	.src0_valid(src0_valid),
	.av_readdata_pre_221(av_readdata_pre_22),
	.av_readdata_pre_23(av_readdata_pre_23),
	.av_readdata_pre_11(av_readdata_pre_11),
	.av_readdata_pre_13(av_readdata_pre_13),
	.av_readdata_pre_161(av_readdata_pre_16),
	.av_readdata_pre_12(av_readdata_pre_12),
	.av_readdata_pre_14(av_readdata_pre_14),
	.av_readdata_pre_15(av_readdata_pre_15),
	.av_readdata_pre_181(av_readdata_pre_18),
	.av_readdata_pre_171(av_readdata_pre_17),
	.av_readdata_pre_10(av_readdata_pre_10),
	.av_readdata_pre_9(av_readdata_pre_9),
	.av_readdata_pre_8(av_readdata_pre_8),
	.av_readdata_pre_211(av_readdata_pre_21),
	.av_readdata_pre_191(av_readdata_pre_19),
	.av_readdata_pre_201(av_readdata_pre_20),
	.av_readdata_pre_81(\avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_82(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[8]~q ),
	.src_data_8(src_data_8),
	.av_readdata_pre_121(\avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_122(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[12]~q ),
	.src_data_12(src_data_12),
	.av_readdata_pre_111(\avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[11]~q ),
	.src_data_11(src_data_11),
	.av_readdata_pre_101(\avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_102(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[10]~q ),
	.src_data_10(src_data_10),
	.av_readdata_pre_91(\avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_92(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[9]~q ),
	.src_data_9(src_data_9),
	.av_readdata_pre_151(\avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_152(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[15]~q ),
	.src_data_15(src_data_15),
	.av_readdata_pre_141(\avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_142(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[14]~q ),
	.src_data_14(src_data_14),
	.av_readdata_pre_131(\avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_132(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[13]~q ),
	.src_data_13(src_data_13),
	.av_readdata_pre_162(\avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[16]~q ),
	.src_data_16(src_data_16),
	.av_readdata_pre_202(\avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[20]~q ),
	.src_data_20(src_data_20),
	.av_readdata_pre_192(\avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[19]~q ),
	.src_data_19(src_data_19),
	.av_readdata_pre_182(\avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[18]~q ),
	.src_data_18(src_data_18),
	.av_readdata_pre_172(\avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[17]~q ),
	.src_data_17(src_data_17),
	.av_readdata_pre_231(\avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[23]~q ),
	.src_data_23(src_data_23),
	.av_readdata_pre_222(\avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[22]~q ),
	.src_data_22(src_data_22),
	.av_readdata_pre_212(\avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[21]~q ),
	.src_data_21(src_data_21));

nios_mcu_nios_mcu_mm_interconnect_0_cmd_demux_001_1 rsp_demux_002(
	.mem_73_0(mem_73_0),
	.mem_55_0(mem_55_0),
	.read_latency_shift_reg_0(read_latency_shift_reg_01),
	.src0_valid(src0_valid),
	.src1_valid(src1_valid));

nios_mcu_altera_merlin_slave_agent avalonslave_0_avalon_slave_0_1_agent(
	.W_alu_result_4(W_alu_result_4),
	.Equal1(Equal1),
	.rst1(rst1),
	.uav_read(\nios_cpu_data_master_translator|uav_read~0_combout ),
	.always2(always2),
	.mem_used_1(\avalonslave_0_avalon_slave_0_1_agent_rsp_fifo|mem_used[1]~q ),
	.m0_read(m0_read),
	.m0_read1(m0_read1));

nios_mcu_altera_avalon_sc_fifo_1 jtag_uart_0_avalon_jtag_slave_agent_rsp_fifo(
	.reset(r_sync_rst),
	.read_latency_shift_reg(read_latency_shift_reg),
	.read_latency_shift_reg_0(read_latency_shift_reg_02),
	.Equal3(Equal3),
	.av_waitrequest(av_waitrequest),
	.mem_used_1(mem_used_13),
	.read_latency_shift_reg1(\jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg~1_combout ),
	.clk(clk_clk));

nios_mcu_altera_merlin_master_agent nios_cpu_data_master_agent(
	.d_write(d_write),
	.write_accepted(write_accepted),
	.d_read(d_read),
	.read_accepted(\nios_cpu_data_master_translator|read_accepted~q ),
	.always2(always2));

nios_mcu_altera_merlin_slave_translator_3 onchip_ram_s1_translator(
	.reset(r_sync_rst),
	.rst1(rst1),
	.F_pc_9(F_pc_9),
	.read_accepted(\nios_cpu_instruction_master_translator|read_accepted~q ),
	.i_read(i_read),
	.read_latency_shift_reg(\onchip_ram_s1_translator|read_latency_shift_reg~0_combout ),
	.Equal0(\router_001|Equal0~0_combout ),
	.read_latency_shift_reg_0(read_latency_shift_reg_05),
	.mem_used_1(\onchip_ram_s1_agent_rsp_fifo|mem_used[1]~q ),
	.read_latency_shift_reg1(\onchip_ram_s1_translator|read_latency_shift_reg~1_combout ),
	.clk(clk_clk));

nios_mcu_altera_merlin_slave_translator_4 onchip_ram_s2_translator(
	.reset(r_sync_rst),
	.read_latency_shift_reg(read_latency_shift_reg),
	.read_latency_shift_reg_0(read_latency_shift_reg_04),
	.src_channel_4(src_channel_4),
	.mem_used_1(mem_used_11),
	.read_latency_shift_reg1(\onchip_ram_s2_translator|read_latency_shift_reg~0_combout ),
	.clk(clk_clk));

nios_mcu_altera_merlin_slave_translator_5 pio_0_s1_translator(
	.W_alu_result_4(W_alu_result_4),
	.reset(r_sync_rst),
	.Equal1(Equal1),
	.mem_used_1(mem_used_1),
	.always0(always0),
	.wait_latency_counter_1(wait_latency_counter_1),
	.wait_latency_counter_0(wait_latency_counter_0),
	.read_latency_shift_reg_0(read_latency_shift_reg_0),
	.read_latency_shift_reg(read_latency_shift_reg),
	.Equal11(\router|Equal1~4_combout ),
	.m0_write(m0_write),
	.wait_latency_counter_11(\pio_0_s1_translator|wait_latency_counter[1]~0_combout ),
	.read_latency_shift_reg1(\pio_0_s1_translator|read_latency_shift_reg~0_combout ),
	.always2(always2),
	.read_latency_shift_reg2(\pio_0_s1_translator|read_latency_shift_reg~1_combout ),
	.av_readdata_pre_0(av_readdata_pre_02),
	.av_readdata_pre_1(av_readdata_pre_112),
	.av_readdata_pre_2(av_readdata_pre_29),
	.av_readdata_pre_3(av_readdata_pre_33),
	.av_readdata_pre_4(av_readdata_pre_43),
	.av_readdata_pre_5(av_readdata_pre_53),
	.av_readdata_pre_6(av_readdata_pre_63),
	.av_readdata_pre_7(av_readdata_pre_73),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_71,readdata_61,readdata_51,readdata_41,readdata_31,readdata_27,readdata_110,readdata_01}),
	.clk(clk_clk));

nios_mcu_altera_merlin_slave_translator_2 nios_cpu_debug_mem_slave_translator(
	.av_readdata({readdata_311,readdata_30,readdata_29,readdata_28,readdata_271,readdata_26,readdata_25,readdata_24,readdata_23,readdata_22,readdata_21,readdata_20,readdata_19,readdata_18,readdata_17,readdata_16,readdata_15,readdata_14,readdata_13,readdata_12,readdata_11,readdata_10,readdata_9,
readdata_8,readdata_7,readdata_6,readdata_5,readdata_4,readdata_3,readdata_2,readdata_1,readdata_0}),
	.reset(r_sync_rst),
	.rst1(rst1),
	.read_latency_shift_reg_0(read_latency_shift_reg_01),
	.write(\nios_cpu_debug_mem_slave_agent_rsp_fifo|write~0_combout ),
	.mem(\nios_cpu_debug_mem_slave_agent_rsp_fifo|mem~1_combout ),
	.WideOr1(WideOr12),
	.av_readdata_pre_0(av_readdata_pre_03),
	.av_readdata_pre_22(av_readdata_pre_22),
	.av_readdata_pre_23(av_readdata_pre_23),
	.av_readdata_pre_24(av_readdata_pre_24),
	.av_readdata_pre_25(av_readdata_pre_25),
	.av_readdata_pre_26(av_readdata_pre_26),
	.av_readdata_pre_11(av_readdata_pre_11),
	.av_readdata_pre_13(av_readdata_pre_13),
	.av_readdata_pre_16(av_readdata_pre_16),
	.av_readdata_pre_12(av_readdata_pre_12),
	.av_readdata_pre_1(av_readdata_pre_1),
	.av_readdata_pre_3(av_readdata_pre_3),
	.av_readdata_pre_2(av_readdata_pre_2),
	.av_readdata_pre_5(av_readdata_pre_5),
	.av_readdata_pre_4(av_readdata_pre_4),
	.av_readdata_pre_14(av_readdata_pre_14),
	.av_readdata_pre_15(av_readdata_pre_15),
	.av_readdata_pre_18(av_readdata_pre_18),
	.av_readdata_pre_17(av_readdata_pre_17),
	.av_readdata_pre_10(av_readdata_pre_10),
	.av_readdata_pre_9(av_readdata_pre_9),
	.av_readdata_pre_8(av_readdata_pre_8),
	.av_readdata_pre_7(av_readdata_pre_7),
	.av_readdata_pre_6(av_readdata_pre_6),
	.av_readdata_pre_21(av_readdata_pre_21),
	.av_readdata_pre_19(av_readdata_pre_19),
	.av_readdata_pre_20(av_readdata_pre_20),
	.av_readdata_pre_27(av_readdata_pre_271),
	.av_readdata_pre_28(av_readdata_pre_281),
	.av_readdata_pre_29(av_readdata_pre_291),
	.av_readdata_pre_30(av_readdata_pre_30),
	.av_readdata_pre_31(av_readdata_pre_311),
	.clk(clk_clk));

nios_mcu_altera_merlin_slave_translator avalonslave_0_avalon_slave_0_1_translator(
	.reset(r_sync_rst),
	.read_latency_shift_reg(read_latency_shift_reg),
	.read_latency_shift_reg_0(read_latency_shift_reg_03),
	.Equal2(Equal2),
	.mem_used_1(\avalonslave_0_avalon_slave_0_1_agent_rsp_fifo|mem_used[1]~q ),
	.Equal21(Equal21),
	.read_latency_shift_reg1(\avalonslave_0_avalon_slave_0_1_translator|read_latency_shift_reg~0_combout ),
	.av_readdata_pre_0(av_readdata_pre_0),
	.av_readdata_pre_1(av_readdata_pre_110),
	.av_readdata_pre_2(av_readdata_pre_27),
	.av_readdata_pre_3(av_readdata_pre_31),
	.av_readdata_pre_4(av_readdata_pre_41),
	.av_readdata_pre_5(av_readdata_pre_51),
	.av_readdata_pre_6(av_readdata_pre_61),
	.av_readdata_pre_7(av_readdata_pre_71),
	.av_readdata_pre_8(\avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[8]~q ),
	.av_readdata({ReadData_31,ReadData_30,ReadData_29,ReadData_28,ReadData_27,ReadData_26,ReadData_25,ReadData_24,ReadData_23,ReadData_22,ReadData_21,ReadData_20,ReadData_19,ReadData_18,ReadData_17,ReadData_16,ReadData_15,ReadData_14,ReadData_13,ReadData_12,ReadData_11,ReadData_10,ReadData_9,
ReadData_8,ReadData_7,ReadData_6,ReadData_5,ReadData_4,ReadData_3,ReadData_2,ReadData_1,ReadData_0}),
	.av_readdata_pre_12(\avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_11(\avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[11]~q ),
	.av_readdata_pre_10(\avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_9(\avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_15(\avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_14(\avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_13(\avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_16(\avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[16]~q ),
	.av_readdata_pre_20(\avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[20]~q ),
	.av_readdata_pre_19(\avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[19]~q ),
	.av_readdata_pre_18(\avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[18]~q ),
	.av_readdata_pre_17(\avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[17]~q ),
	.av_readdata_pre_23(\avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[23]~q ),
	.av_readdata_pre_22(\avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[22]~q ),
	.av_readdata_pre_21(\avalonslave_0_avalon_slave_0_1_translator|av_readdata_pre[21]~q ),
	.av_readdata_pre_24(av_readdata_pre_241),
	.av_readdata_pre_31(av_readdata_pre_312),
	.av_readdata_pre_30(av_readdata_pre_301),
	.av_readdata_pre_29(av_readdata_pre_292),
	.av_readdata_pre_28(av_readdata_pre_282),
	.av_readdata_pre_27(av_readdata_pre_272),
	.av_readdata_pre_26(av_readdata_pre_261),
	.av_readdata_pre_25(av_readdata_pre_251),
	.clk(clk_clk));

nios_mcu_altera_merlin_slave_translator_1 jtag_uart_0_avalon_jtag_slave_translator(
	.av_readdata_pre_16(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[16]~q ),
	.av_readdata_pre_20(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[20]~q ),
	.av_readdata_pre_19(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[19]~q ),
	.av_readdata_pre_18(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[18]~q ),
	.av_readdata_pre_17(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[17]~q ),
	.av_readdata_pre_22(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[22]~q ),
	.av_readdata_pre_21(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[21]~q ),
	.reset(r_sync_rst),
	.rst1(rst1),
	.d_read(d_read),
	.read_accepted(\nios_cpu_data_master_translator|read_accepted~q ),
	.read_latency_shift_reg(read_latency_shift_reg),
	.read_latency_shift_reg_0(read_latency_shift_reg_02),
	.Equal3(Equal3),
	.av_waitrequest(av_waitrequest),
	.mem_used_1(mem_used_13),
	.read_latency_shift_reg1(\jtag_uart_0_avalon_jtag_slave_translator|read_latency_shift_reg~1_combout ),
	.av_readdata_pre_0(av_readdata_pre_01),
	.av_readdata_pre_1(av_readdata_pre_111),
	.av_readdata_pre_2(av_readdata_pre_28),
	.av_readdata_pre_3(av_readdata_pre_32),
	.av_readdata_pre_4(av_readdata_pre_42),
	.av_readdata_pre_5(av_readdata_pre_52),
	.av_readdata_pre_6(av_readdata_pre_62),
	.av_readdata_pre_7(av_readdata_pre_72),
	.b_full(b_full),
	.av_readdata_pre_8(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[8]~q ),
	.read_0(read_0),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,rvalid,woverflow,gnd,b_non_empty,gnd,ac,av_readdata_9,av_readdata_8,av_readdata_7,av_readdata_6,av_readdata_5,av_readdata_4,av_readdata_3,av_readdata_2,av_readdata_1,av_readdata_0}),
	.av_readdata_pre_12(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_10(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_9(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_15(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_14(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_13(\jtag_uart_0_avalon_jtag_slave_translator|av_readdata_pre[13]~q ),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_31(counter_reg_bit_31),
	.counter_reg_bit_01(counter_reg_bit_01),
	.counter_reg_bit_21(counter_reg_bit_21),
	.counter_reg_bit_11(counter_reg_bit_11),
	.b_full1(b_full1),
	.counter_reg_bit_51(counter_reg_bit_51),
	.counter_reg_bit_41(counter_reg_bit_41),
	.clk(clk_clk));

nios_mcu_altera_merlin_master_translator_1 nios_cpu_instruction_master_translator(
	.reset(r_sync_rst),
	.rst1(rst1),
	.write(\nios_cpu_debug_mem_slave_agent_rsp_fifo|write~0_combout ),
	.saved_grant_1(\cmd_mux_002|saved_grant[1]~q ),
	.read_accepted1(\nios_cpu_instruction_master_translator|read_accepted~q ),
	.i_read(i_read),
	.read_latency_shift_reg_0(read_latency_shift_reg_05),
	.src1_valid(src1_valid),
	.Equal0(\router_001|Equal0~1_combout ),
	.mem_used_1(\onchip_ram_s1_agent_rsp_fifo|mem_used[1]~q ),
	.clk(clk_clk));

nios_mcu_altera_merlin_master_translator nios_cpu_data_master_translator(
	.reset(r_sync_rst),
	.rst1(rst1),
	.d_write(d_write),
	.write_accepted1(write_accepted),
	.d_read(d_read),
	.read_accepted1(\nios_cpu_data_master_translator|read_accepted~q ),
	.WideOr1(WideOr11),
	.sink_ready(\cmd_demux|sink_ready~0_combout ),
	.WideOr0(\cmd_demux|WideOr0~0_combout ),
	.read_latency_shift_reg(\pio_0_s1_translator|read_latency_shift_reg~0_combout ),
	.uav_read(\nios_cpu_data_master_translator|uav_read~0_combout ),
	.always2(always2),
	.sink_ready1(\cmd_demux|sink_ready~2_combout ),
	.av_waitrequest(nios_cpu_data_master_waitrequest),
	.WideOr01(\cmd_demux|WideOr0~1_combout ),
	.clk(clk_clk));

endmodule

module nios_mcu_altera_avalon_sc_fifo (
	reset,
	rst1,
	read_latency_shift_reg_0,
	Equal2,
	uav_read,
	mem_used_1,
	Equal21,
	read_latency_shift_reg,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	rst1;
input 	read_latency_shift_reg_0;
input 	Equal2;
input 	uav_read;
output 	mem_used_1;
input 	Equal21;
input 	read_latency_shift_reg;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~2_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem_used[1]~1_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cycloneive_lcell_comb \mem_used[0]~2 (
	.dataa(read_latency_shift_reg),
	.datab(\mem_used[0]~q ),
	.datac(mem_used_1),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[0]~2_combout ),
	.cout());
defparam \mem_used[0]~2 .lut_mask = 16'hFEFF;
defparam \mem_used[0]~2 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cycloneive_lcell_comb \mem_used[1]~0 (
	.dataa(rst1),
	.datab(uav_read),
	.datac(Equal2),
	.datad(Equal21),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hFEFF;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~1 (
	.dataa(mem_used_1),
	.datab(read_latency_shift_reg_0),
	.datac(\mem_used[0]~q ),
	.datad(\mem_used[1]~0_combout ),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hBFB3;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

endmodule

module nios_mcu_altera_avalon_sc_fifo_1 (
	reset,
	read_latency_shift_reg,
	read_latency_shift_reg_0,
	Equal3,
	av_waitrequest,
	mem_used_1,
	read_latency_shift_reg1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	read_latency_shift_reg;
input 	read_latency_shift_reg_0;
input 	Equal3;
input 	av_waitrequest;
output 	mem_used_1;
input 	read_latency_shift_reg1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~2_combout ;
wire \mem_used[0]~3_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem_used[1]~1_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cycloneive_lcell_comb \mem_used[0]~2 (
	.dataa(Equal3),
	.datab(read_latency_shift_reg),
	.datac(av_waitrequest),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_used[0]~2_combout ),
	.cout());
defparam \mem_used[0]~2 .lut_mask = 16'hFEFE;
defparam \mem_used[0]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~3 (
	.dataa(\mem_used[0]~q ),
	.datab(mem_used_1),
	.datac(read_latency_shift_reg_0),
	.datad(\mem_used[0]~2_combout ),
	.cin(gnd),
	.combout(\mem_used[0]~3_combout ),
	.cout());
defparam \mem_used[0]~3 .lut_mask = 16'hBF8F;
defparam \mem_used[0]~3 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cycloneive_lcell_comb \mem_used[1]~0 (
	.dataa(Equal3),
	.datab(\mem_used[0]~q ),
	.datac(read_latency_shift_reg1),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hFEFF;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~1 (
	.dataa(\mem_used[1]~0_combout ),
	.datab(mem_used_1),
	.datac(read_latency_shift_reg_0),
	.datad(\mem_used[0]~q ),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hEFFF;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

endmodule

module nios_mcu_altera_avalon_sc_fifo_2 (
	reset,
	mem_73_0,
	mem_55_0,
	read_latency_shift_reg_0,
	waitrequest,
	mem_used_1,
	write,
	saved_grant_1,
	rf_source_valid,
	read_accepted,
	i_read,
	mem,
	WideOr1,
	rf_source_valid1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
output 	mem_73_0;
output 	mem_55_0;
input 	read_latency_shift_reg_0;
input 	waitrequest;
output 	mem_used_1;
output 	write;
input 	saved_grant_1;
input 	rf_source_valid;
input 	read_accepted;
input 	i_read;
output 	mem;
input 	WideOr1;
input 	rf_source_valid1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem[1][73]~q ;
wire \mem~0_combout ;
wire \mem_used[0]~3_combout ;
wire \mem_used[0]~4_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem[1][55]~q ;
wire \mem~2_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~2_combout ;


dffeas \mem[0][73] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_73_0),
	.prn(vcc));
defparam \mem[0][73] .is_wysiwyg = "true";
defparam \mem[0][73] .power_up = "low";

dffeas \mem[0][55] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_55_0),
	.prn(vcc));
defparam \mem[0][55] .is_wysiwyg = "true";
defparam \mem[0][55] .power_up = "low";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cycloneive_lcell_comb \write~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(waitrequest),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(write),
	.cout());
defparam \write~0 .lut_mask = 16'h0FFF;
defparam \write~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem~1 (
	.dataa(rf_source_valid),
	.datab(saved_grant_1),
	.datac(read_accepted),
	.datad(i_read),
	.cin(gnd),
	.combout(mem),
	.cout());
defparam \mem~1 .lut_mask = 16'hEFFF;
defparam \mem~1 .sum_lutc_input = "datac";

dffeas \mem[1][73] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][73]~q ),
	.prn(vcc));
defparam \mem[1][73] .is_wysiwyg = "true";
defparam \mem[1][73] .power_up = "low";

cycloneive_lcell_comb \mem~0 (
	.dataa(\mem[1][73]~q ),
	.datab(saved_grant_1),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~0_combout ),
	.cout());
defparam \mem~0 .lut_mask = 16'hAACC;
defparam \mem~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~3 (
	.dataa(\mem_used[0]~q ),
	.datab(mem_used_1),
	.datac(gnd),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[0]~3_combout ),
	.cout());
defparam \mem_used[0]~3 .lut_mask = 16'hEEFF;
defparam \mem_used[0]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[0]~4 (
	.dataa(\mem_used[0]~3_combout ),
	.datab(write),
	.datac(WideOr1),
	.datad(mem),
	.cin(gnd),
	.combout(\mem_used[0]~4_combout ),
	.cout());
defparam \mem_used[0]~4 .lut_mask = 16'hFFFE;
defparam \mem_used[0]~4 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cycloneive_lcell_comb \mem_used[1]~0 (
	.dataa(\mem_used[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hFF55;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

dffeas \mem[1][55] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][55]~q ),
	.prn(vcc));
defparam \mem[1][55] .is_wysiwyg = "true";
defparam \mem[1][55] .power_up = "low";

cycloneive_lcell_comb \mem~2 (
	.dataa(\mem[1][55]~q ),
	.datab(mem),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~2_combout ),
	.cout());
defparam \mem~2 .lut_mask = 16'hAACC;
defparam \mem~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~1 (
	.dataa(mem_used_1),
	.datab(gnd),
	.datac(read_latency_shift_reg_0),
	.datad(\mem_used[0]~q ),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hAFFF;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~2 (
	.dataa(\mem_used[1]~1_combout ),
	.datab(rf_source_valid1),
	.datac(\mem_used[1]~0_combout ),
	.datad(waitrequest),
	.cin(gnd),
	.combout(\mem_used[1]~2_combout ),
	.cout());
defparam \mem_used[1]~2 .lut_mask = 16'hEFFF;
defparam \mem_used[1]~2 .sum_lutc_input = "datac";

endmodule

module nios_mcu_altera_avalon_sc_fifo_3 (
	reset,
	read_latency_shift_reg,
	read_latency_shift_reg_0,
	Equal0,
	mem_used_1,
	read_latency_shift_reg1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	read_latency_shift_reg;
input 	read_latency_shift_reg_0;
input 	Equal0;
output 	mem_used_1;
input 	read_latency_shift_reg1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~2_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem_used[1]~1_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cycloneive_lcell_comb \mem_used[0]~2 (
	.dataa(read_latency_shift_reg1),
	.datab(\mem_used[0]~q ),
	.datac(mem_used_1),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[0]~2_combout ),
	.cout());
defparam \mem_used[0]~2 .lut_mask = 16'hFEFF;
defparam \mem_used[0]~2 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cycloneive_lcell_comb \mem_used[1]~0 (
	.dataa(read_latency_shift_reg),
	.datab(\mem_used[0]~q ),
	.datac(Equal0),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hEFFF;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~1 (
	.dataa(\mem_used[1]~0_combout ),
	.datab(mem_used_1),
	.datac(read_latency_shift_reg_0),
	.datad(\mem_used[0]~q ),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hEFFF;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

endmodule

module nios_mcu_altera_avalon_sc_fifo_4 (
	reset,
	read_latency_shift_reg,
	read_latency_shift_reg_0,
	src_channel_4,
	mem_used_1,
	read_latency_shift_reg1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	read_latency_shift_reg;
input 	read_latency_shift_reg_0;
input 	src_channel_4;
output 	mem_used_1;
input 	read_latency_shift_reg1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~2_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem_used[1]~1_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cycloneive_lcell_comb \mem_used[0]~2 (
	.dataa(read_latency_shift_reg1),
	.datab(\mem_used[0]~q ),
	.datac(mem_used_1),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[0]~2_combout ),
	.cout());
defparam \mem_used[0]~2 .lut_mask = 16'hFEFF;
defparam \mem_used[0]~2 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cycloneive_lcell_comb \mem_used[1]~0 (
	.dataa(read_latency_shift_reg),
	.datab(src_channel_4),
	.datac(\mem_used[0]~q ),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hFEFF;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~1 (
	.dataa(\mem_used[1]~0_combout ),
	.datab(mem_used_1),
	.datac(read_latency_shift_reg_0),
	.datad(\mem_used[0]~q ),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hEFFF;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

endmodule

module nios_mcu_altera_avalon_sc_fifo_5 (
	W_alu_result_4,
	reset,
	Equal1,
	mem_used_1,
	read_latency_shift_reg_0,
	read_latency_shift_reg,
	wait_latency_counter_1,
	read_latency_shift_reg1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_4;
input 	reset;
input 	Equal1;
output 	mem_used_1;
input 	read_latency_shift_reg_0;
input 	read_latency_shift_reg;
input 	wait_latency_counter_1;
input 	read_latency_shift_reg1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~3_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~4_combout ;
wire \mem_used[1]~2_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cycloneive_lcell_comb \mem_used[0]~3 (
	.dataa(read_latency_shift_reg1),
	.datab(\mem_used[0]~q ),
	.datac(mem_used_1),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[0]~3_combout ),
	.cout());
defparam \mem_used[0]~3 .lut_mask = 16'hFEFF;
defparam \mem_used[0]~3 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cycloneive_lcell_comb \mem_used[1]~4 (
	.dataa(Equal1),
	.datab(W_alu_result_4),
	.datac(read_latency_shift_reg),
	.datad(wait_latency_counter_1),
	.cin(gnd),
	.combout(\mem_used[1]~4_combout ),
	.cout());
defparam \mem_used[1]~4 .lut_mask = 16'hFFFB;
defparam \mem_used[1]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[1]~2 (
	.dataa(mem_used_1),
	.datab(read_latency_shift_reg_0),
	.datac(\mem_used[0]~q ),
	.datad(\mem_used[1]~4_combout ),
	.cin(gnd),
	.combout(\mem_used[1]~2_combout ),
	.cout());
defparam \mem_used[1]~2 .lut_mask = 16'hBFB3;
defparam \mem_used[1]~2 .sum_lutc_input = "datac";

endmodule

module nios_mcu_altera_merlin_master_agent (
	d_write,
	write_accepted,
	d_read,
	read_accepted,
	always2)/* synthesis synthesis_greybox=1 */;
input 	d_write;
input 	write_accepted;
input 	d_read;
input 	read_accepted;
output 	always2;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \always2~0 (
	.dataa(d_write),
	.datab(d_read),
	.datac(write_accepted),
	.datad(read_accepted),
	.cin(gnd),
	.combout(always2),
	.cout());
defparam \always2~0 .lut_mask = 16'hEFFF;
defparam \always2~0 .sum_lutc_input = "datac";

endmodule

module nios_mcu_altera_merlin_master_translator (
	reset,
	rst1,
	d_write,
	write_accepted1,
	d_read,
	read_accepted1,
	WideOr1,
	sink_ready,
	WideOr0,
	read_latency_shift_reg,
	uav_read,
	always2,
	sink_ready1,
	av_waitrequest,
	WideOr01,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	rst1;
input 	d_write;
output 	write_accepted1;
input 	d_read;
output 	read_accepted1;
input 	WideOr1;
input 	sink_ready;
input 	WideOr0;
input 	read_latency_shift_reg;
output 	uav_read;
input 	always2;
input 	sink_ready1;
output 	av_waitrequest;
input 	WideOr01;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_accepted~0_combout ;
wire \write_accepted~0_combout ;
wire \read_accepted~1_combout ;
wire \end_begintransfer~0_combout ;
wire \end_begintransfer~q ;
wire \av_waitrequest~0_combout ;
wire \av_waitrequest~1_combout ;


dffeas write_accepted(
	.clk(clk),
	.d(\write_accepted~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(write_accepted1),
	.prn(vcc));
defparam write_accepted.is_wysiwyg = "true";
defparam write_accepted.power_up = "low";

dffeas read_accepted(
	.clk(clk),
	.d(\read_accepted~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_accepted1),
	.prn(vcc));
defparam read_accepted.is_wysiwyg = "true";
defparam read_accepted.power_up = "low";

cycloneive_lcell_comb \uav_read~0 (
	.dataa(d_read),
	.datab(gnd),
	.datac(gnd),
	.datad(read_accepted1),
	.cin(gnd),
	.combout(uav_read),
	.cout());
defparam \uav_read~0 .lut_mask = 16'hAAFF;
defparam \uav_read~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_waitrequest~2 (
	.dataa(d_read),
	.datab(WideOr1),
	.datac(d_write),
	.datad(\av_waitrequest~1_combout ),
	.cin(gnd),
	.combout(av_waitrequest),
	.cout());
defparam \av_waitrequest~2 .lut_mask = 16'h8DFF;
defparam \av_waitrequest~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_accepted~0 (
	.dataa(rst1),
	.datab(sink_ready1),
	.datac(read_latency_shift_reg),
	.datad(WideOr01),
	.cin(gnd),
	.combout(\read_accepted~0_combout ),
	.cout());
defparam \read_accepted~0 .lut_mask = 16'hFFFE;
defparam \read_accepted~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \write_accepted~0 (
	.dataa(av_waitrequest),
	.datab(write_accepted1),
	.datac(d_write),
	.datad(\read_accepted~0_combout ),
	.cin(gnd),
	.combout(\write_accepted~0_combout ),
	.cout());
defparam \write_accepted~0 .lut_mask = 16'hFFFE;
defparam \write_accepted~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_accepted~1 (
	.dataa(WideOr1),
	.datab(read_accepted1),
	.datac(d_read),
	.datad(\read_accepted~0_combout ),
	.cin(gnd),
	.combout(\read_accepted~1_combout ),
	.cout());
defparam \read_accepted~1 .lut_mask = 16'hFFFE;
defparam \read_accepted~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \end_begintransfer~0 (
	.dataa(always2),
	.datab(\end_begintransfer~q ),
	.datac(gnd),
	.datad(\read_accepted~0_combout ),
	.cin(gnd),
	.combout(\end_begintransfer~0_combout ),
	.cout());
defparam \end_begintransfer~0 .lut_mask = 16'hEEFF;
defparam \end_begintransfer~0 .sum_lutc_input = "datac";

dffeas end_begintransfer(
	.clk(clk),
	.d(\end_begintransfer~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\end_begintransfer~q ),
	.prn(vcc));
defparam end_begintransfer.is_wysiwyg = "true";
defparam end_begintransfer.power_up = "low";

cycloneive_lcell_comb \av_waitrequest~0 (
	.dataa(sink_ready),
	.datab(WideOr0),
	.datac(read_latency_shift_reg),
	.datad(sink_ready1),
	.cin(gnd),
	.combout(\av_waitrequest~0_combout ),
	.cout());
defparam \av_waitrequest~0 .lut_mask = 16'hFFFE;
defparam \av_waitrequest~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_waitrequest~1 (
	.dataa(rst1),
	.datab(\end_begintransfer~q ),
	.datac(write_accepted1),
	.datad(\av_waitrequest~0_combout ),
	.cin(gnd),
	.combout(\av_waitrequest~1_combout ),
	.cout());
defparam \av_waitrequest~1 .lut_mask = 16'hFFFE;
defparam \av_waitrequest~1 .sum_lutc_input = "datac";

endmodule

module nios_mcu_altera_merlin_master_translator_1 (
	reset,
	rst1,
	write,
	saved_grant_1,
	read_accepted1,
	i_read,
	read_latency_shift_reg_0,
	src1_valid,
	Equal0,
	mem_used_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	rst1;
input 	write;
input 	saved_grant_1;
output 	read_accepted1;
input 	i_read;
input 	read_latency_shift_reg_0;
input 	src1_valid;
input 	Equal0;
input 	mem_used_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_accepted~0_combout ;
wire \read_accepted~1_combout ;
wire \read_accepted~2_combout ;


dffeas read_accepted(
	.clk(clk),
	.d(\read_accepted~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_accepted1),
	.prn(vcc));
defparam read_accepted.is_wysiwyg = "true";
defparam read_accepted.power_up = "low";

cycloneive_lcell_comb \read_accepted~0 (
	.dataa(write),
	.datab(saved_grant_1),
	.datac(Equal0),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\read_accepted~0_combout ),
	.cout());
defparam \read_accepted~0 .lut_mask = 16'hACFF;
defparam \read_accepted~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_accepted~1 (
	.dataa(read_accepted1),
	.datab(rst1),
	.datac(\read_accepted~0_combout ),
	.datad(i_read),
	.cin(gnd),
	.combout(\read_accepted~1_combout ),
	.cout());
defparam \read_accepted~1 .lut_mask = 16'hFEFF;
defparam \read_accepted~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_accepted~2 (
	.dataa(\read_accepted~1_combout ),
	.datab(gnd),
	.datac(src1_valid),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\read_accepted~2_combout ),
	.cout());
defparam \read_accepted~2 .lut_mask = 16'hAFFF;
defparam \read_accepted~2 .sum_lutc_input = "datac";

endmodule

module nios_mcu_altera_merlin_slave_agent (
	W_alu_result_4,
	Equal1,
	rst1,
	uav_read,
	always2,
	mem_used_1,
	m0_read,
	m0_read1)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_4;
input 	Equal1;
input 	rst1;
input 	uav_read;
input 	always2;
input 	mem_used_1;
output 	m0_read;
output 	m0_read1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \m0_read~0 (
	.dataa(rst1),
	.datab(always2),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(m0_read),
	.cout());
defparam \m0_read~0 .lut_mask = 16'hEEFF;
defparam \m0_read~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \m0_read~1 (
	.dataa(W_alu_result_4),
	.datab(Equal1),
	.datac(uav_read),
	.datad(m0_read),
	.cin(gnd),
	.combout(m0_read1),
	.cout());
defparam \m0_read~1 .lut_mask = 16'hFFFE;
defparam \m0_read~1 .sum_lutc_input = "datac";

endmodule

module nios_mcu_altera_merlin_slave_agent_2 (
	d_read,
	read_accepted,
	saved_grant_0,
	rf_source_valid,
	mem,
	WideOr1,
	rf_source_valid1)/* synthesis synthesis_greybox=1 */;
input 	d_read;
input 	read_accepted;
input 	saved_grant_0;
output 	rf_source_valid;
input 	mem;
input 	WideOr1;
output 	rf_source_valid1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \rf_source_valid~0 (
	.dataa(d_read),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(read_accepted),
	.cin(gnd),
	.combout(rf_source_valid),
	.cout());
defparam \rf_source_valid~0 .lut_mask = 16'hEEFF;
defparam \rf_source_valid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rf_source_valid~1 (
	.dataa(WideOr1),
	.datab(mem),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(rf_source_valid1),
	.cout());
defparam \rf_source_valid~1 .lut_mask = 16'hEEEE;
defparam \rf_source_valid~1 .sum_lutc_input = "datac";

endmodule

module nios_mcu_altera_merlin_slave_agent_5 (
	d_write,
	write_accepted,
	m0_write)/* synthesis synthesis_greybox=1 */;
input 	d_write;
input 	write_accepted;
output 	m0_write;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \m0_write~0 (
	.dataa(d_write),
	.datab(gnd),
	.datac(gnd),
	.datad(write_accepted),
	.cin(gnd),
	.combout(m0_write),
	.cout());
defparam \m0_write~0 .lut_mask = 16'hAAFF;
defparam \m0_write~0 .sum_lutc_input = "datac";

endmodule

module nios_mcu_altera_merlin_slave_translator (
	reset,
	read_latency_shift_reg,
	read_latency_shift_reg_0,
	Equal2,
	mem_used_1,
	Equal21,
	read_latency_shift_reg1,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata_pre_8,
	av_readdata,
	av_readdata_pre_12,
	av_readdata_pre_11,
	av_readdata_pre_10,
	av_readdata_pre_9,
	av_readdata_pre_15,
	av_readdata_pre_14,
	av_readdata_pre_13,
	av_readdata_pre_16,
	av_readdata_pre_20,
	av_readdata_pre_19,
	av_readdata_pre_18,
	av_readdata_pre_17,
	av_readdata_pre_23,
	av_readdata_pre_22,
	av_readdata_pre_21,
	av_readdata_pre_24,
	av_readdata_pre_31,
	av_readdata_pre_30,
	av_readdata_pre_29,
	av_readdata_pre_28,
	av_readdata_pre_27,
	av_readdata_pre_26,
	av_readdata_pre_25,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	read_latency_shift_reg;
output 	read_latency_shift_reg_0;
input 	Equal2;
input 	mem_used_1;
input 	Equal21;
output 	read_latency_shift_reg1;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
output 	av_readdata_pre_8;
input 	[31:0] av_readdata;
output 	av_readdata_pre_12;
output 	av_readdata_pre_11;
output 	av_readdata_pre_10;
output 	av_readdata_pre_9;
output 	av_readdata_pre_15;
output 	av_readdata_pre_14;
output 	av_readdata_pre_13;
output 	av_readdata_pre_16;
output 	av_readdata_pre_20;
output 	av_readdata_pre_19;
output 	av_readdata_pre_18;
output 	av_readdata_pre_17;
output 	av_readdata_pre_23;
output 	av_readdata_pre_22;
output 	av_readdata_pre_21;
output 	av_readdata_pre_24;
output 	av_readdata_pre_31;
output 	av_readdata_pre_30;
output 	av_readdata_pre_29;
output 	av_readdata_pre_28;
output 	av_readdata_pre_27;
output 	av_readdata_pre_26;
output 	av_readdata_pre_25;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(read_latency_shift_reg1),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cycloneive_lcell_comb \read_latency_shift_reg~0 (
	.dataa(read_latency_shift_reg),
	.datab(Equal2),
	.datac(mem_used_1),
	.datad(Equal21),
	.cin(gnd),
	.combout(read_latency_shift_reg1),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hEFFF;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[12] (
	.clk(clk),
	.d(av_readdata[12]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_12),
	.prn(vcc));
defparam \av_readdata_pre[12] .is_wysiwyg = "true";
defparam \av_readdata_pre[12] .power_up = "low";

dffeas \av_readdata_pre[11] (
	.clk(clk),
	.d(av_readdata[11]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_11),
	.prn(vcc));
defparam \av_readdata_pre[11] .is_wysiwyg = "true";
defparam \av_readdata_pre[11] .power_up = "low";

dffeas \av_readdata_pre[10] (
	.clk(clk),
	.d(av_readdata[10]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_10),
	.prn(vcc));
defparam \av_readdata_pre[10] .is_wysiwyg = "true";
defparam \av_readdata_pre[10] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[15] (
	.clk(clk),
	.d(av_readdata[15]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_15),
	.prn(vcc));
defparam \av_readdata_pre[15] .is_wysiwyg = "true";
defparam \av_readdata_pre[15] .power_up = "low";

dffeas \av_readdata_pre[14] (
	.clk(clk),
	.d(av_readdata[14]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_14),
	.prn(vcc));
defparam \av_readdata_pre[14] .is_wysiwyg = "true";
defparam \av_readdata_pre[14] .power_up = "low";

dffeas \av_readdata_pre[13] (
	.clk(clk),
	.d(av_readdata[13]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_13),
	.prn(vcc));
defparam \av_readdata_pre[13] .is_wysiwyg = "true";
defparam \av_readdata_pre[13] .power_up = "low";

dffeas \av_readdata_pre[16] (
	.clk(clk),
	.d(av_readdata[16]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_16),
	.prn(vcc));
defparam \av_readdata_pre[16] .is_wysiwyg = "true";
defparam \av_readdata_pre[16] .power_up = "low";

dffeas \av_readdata_pre[20] (
	.clk(clk),
	.d(av_readdata[20]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_20),
	.prn(vcc));
defparam \av_readdata_pre[20] .is_wysiwyg = "true";
defparam \av_readdata_pre[20] .power_up = "low";

dffeas \av_readdata_pre[19] (
	.clk(clk),
	.d(av_readdata[19]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_19),
	.prn(vcc));
defparam \av_readdata_pre[19] .is_wysiwyg = "true";
defparam \av_readdata_pre[19] .power_up = "low";

dffeas \av_readdata_pre[18] (
	.clk(clk),
	.d(av_readdata[18]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_18),
	.prn(vcc));
defparam \av_readdata_pre[18] .is_wysiwyg = "true";
defparam \av_readdata_pre[18] .power_up = "low";

dffeas \av_readdata_pre[17] (
	.clk(clk),
	.d(av_readdata[17]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_17),
	.prn(vcc));
defparam \av_readdata_pre[17] .is_wysiwyg = "true";
defparam \av_readdata_pre[17] .power_up = "low";

dffeas \av_readdata_pre[23] (
	.clk(clk),
	.d(av_readdata[23]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_23),
	.prn(vcc));
defparam \av_readdata_pre[23] .is_wysiwyg = "true";
defparam \av_readdata_pre[23] .power_up = "low";

dffeas \av_readdata_pre[22] (
	.clk(clk),
	.d(av_readdata[22]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_22),
	.prn(vcc));
defparam \av_readdata_pre[22] .is_wysiwyg = "true";
defparam \av_readdata_pre[22] .power_up = "low";

dffeas \av_readdata_pre[21] (
	.clk(clk),
	.d(av_readdata[21]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_21),
	.prn(vcc));
defparam \av_readdata_pre[21] .is_wysiwyg = "true";
defparam \av_readdata_pre[21] .power_up = "low";

dffeas \av_readdata_pre[24] (
	.clk(clk),
	.d(av_readdata[24]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_24),
	.prn(vcc));
defparam \av_readdata_pre[24] .is_wysiwyg = "true";
defparam \av_readdata_pre[24] .power_up = "low";

dffeas \av_readdata_pre[31] (
	.clk(clk),
	.d(av_readdata[31]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_31),
	.prn(vcc));
defparam \av_readdata_pre[31] .is_wysiwyg = "true";
defparam \av_readdata_pre[31] .power_up = "low";

dffeas \av_readdata_pre[30] (
	.clk(clk),
	.d(av_readdata[30]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_30),
	.prn(vcc));
defparam \av_readdata_pre[30] .is_wysiwyg = "true";
defparam \av_readdata_pre[30] .power_up = "low";

dffeas \av_readdata_pre[29] (
	.clk(clk),
	.d(av_readdata[29]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_29),
	.prn(vcc));
defparam \av_readdata_pre[29] .is_wysiwyg = "true";
defparam \av_readdata_pre[29] .power_up = "low";

dffeas \av_readdata_pre[28] (
	.clk(clk),
	.d(av_readdata[28]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_28),
	.prn(vcc));
defparam \av_readdata_pre[28] .is_wysiwyg = "true";
defparam \av_readdata_pre[28] .power_up = "low";

dffeas \av_readdata_pre[27] (
	.clk(clk),
	.d(av_readdata[27]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_27),
	.prn(vcc));
defparam \av_readdata_pre[27] .is_wysiwyg = "true";
defparam \av_readdata_pre[27] .power_up = "low";

dffeas \av_readdata_pre[26] (
	.clk(clk),
	.d(av_readdata[26]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_26),
	.prn(vcc));
defparam \av_readdata_pre[26] .is_wysiwyg = "true";
defparam \av_readdata_pre[26] .power_up = "low";

dffeas \av_readdata_pre[25] (
	.clk(clk),
	.d(av_readdata[25]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_25),
	.prn(vcc));
defparam \av_readdata_pre[25] .is_wysiwyg = "true";
defparam \av_readdata_pre[25] .power_up = "low";

endmodule

module nios_mcu_altera_merlin_slave_translator_1 (
	av_readdata_pre_16,
	av_readdata_pre_20,
	av_readdata_pre_19,
	av_readdata_pre_18,
	av_readdata_pre_17,
	av_readdata_pre_22,
	av_readdata_pre_21,
	reset,
	rst1,
	d_read,
	read_accepted,
	read_latency_shift_reg,
	read_latency_shift_reg_0,
	Equal3,
	av_waitrequest,
	mem_used_1,
	read_latency_shift_reg1,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	b_full,
	av_readdata_pre_8,
	read_0,
	av_readdata,
	av_readdata_pre_12,
	av_readdata_pre_10,
	av_readdata_pre_9,
	av_readdata_pre_15,
	av_readdata_pre_14,
	av_readdata_pre_13,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_31,
	counter_reg_bit_01,
	counter_reg_bit_21,
	counter_reg_bit_11,
	b_full1,
	counter_reg_bit_51,
	counter_reg_bit_41,
	clk)/* synthesis synthesis_greybox=1 */;
output 	av_readdata_pre_16;
output 	av_readdata_pre_20;
output 	av_readdata_pre_19;
output 	av_readdata_pre_18;
output 	av_readdata_pre_17;
output 	av_readdata_pre_22;
output 	av_readdata_pre_21;
input 	reset;
input 	rst1;
input 	d_read;
input 	read_accepted;
output 	read_latency_shift_reg;
output 	read_latency_shift_reg_0;
input 	Equal3;
input 	av_waitrequest;
input 	mem_used_1;
output 	read_latency_shift_reg1;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
input 	b_full;
output 	av_readdata_pre_8;
input 	read_0;
input 	[31:0] av_readdata;
output 	av_readdata_pre_12;
output 	av_readdata_pre_10;
output 	av_readdata_pre_9;
output 	av_readdata_pre_15;
output 	av_readdata_pre_14;
output 	av_readdata_pre_13;
input 	counter_reg_bit_5;
input 	counter_reg_bit_4;
input 	counter_reg_bit_3;
input 	counter_reg_bit_2;
input 	counter_reg_bit_1;
input 	counter_reg_bit_0;
input 	counter_reg_bit_31;
input 	counter_reg_bit_01;
input 	counter_reg_bit_21;
input 	counter_reg_bit_11;
input 	b_full1;
input 	counter_reg_bit_51;
input 	counter_reg_bit_41;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \av_readdata_pre[16]~7_combout ;
wire \av_readdata_pre[16]~8 ;
wire \av_readdata_pre[17]~10 ;
wire \av_readdata_pre[18]~12 ;
wire \av_readdata_pre[19]~14 ;
wire \av_readdata_pre[20]~15_combout ;
wire \av_readdata_pre[19]~13_combout ;
wire \av_readdata_pre[18]~11_combout ;
wire \av_readdata_pre[17]~9_combout ;
wire \av_readdata_pre[20]~16 ;
wire \av_readdata_pre[21]~18 ;
wire \av_readdata_pre[22]~19_combout ;
wire \av_readdata_pre[21]~17_combout ;
wire \read_latency_shift_reg~2_combout ;
wire \av_readdata_pre[13]~21_combout ;


dffeas \av_readdata_pre[16] (
	.clk(clk),
	.d(\av_readdata_pre[16]~7_combout ),
	.asdata(counter_reg_bit_0),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_16),
	.prn(vcc));
defparam \av_readdata_pre[16] .is_wysiwyg = "true";
defparam \av_readdata_pre[16] .power_up = "low";

dffeas \av_readdata_pre[20] (
	.clk(clk),
	.d(\av_readdata_pre[20]~15_combout ),
	.asdata(counter_reg_bit_4),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_20),
	.prn(vcc));
defparam \av_readdata_pre[20] .is_wysiwyg = "true";
defparam \av_readdata_pre[20] .power_up = "low";

dffeas \av_readdata_pre[19] (
	.clk(clk),
	.d(\av_readdata_pre[19]~13_combout ),
	.asdata(counter_reg_bit_3),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_19),
	.prn(vcc));
defparam \av_readdata_pre[19] .is_wysiwyg = "true";
defparam \av_readdata_pre[19] .power_up = "low";

dffeas \av_readdata_pre[18] (
	.clk(clk),
	.d(\av_readdata_pre[18]~11_combout ),
	.asdata(counter_reg_bit_2),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_18),
	.prn(vcc));
defparam \av_readdata_pre[18] .is_wysiwyg = "true";
defparam \av_readdata_pre[18] .power_up = "low";

dffeas \av_readdata_pre[17] (
	.clk(clk),
	.d(\av_readdata_pre[17]~9_combout ),
	.asdata(counter_reg_bit_1),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_17),
	.prn(vcc));
defparam \av_readdata_pre[17] .is_wysiwyg = "true";
defparam \av_readdata_pre[17] .power_up = "low";

dffeas \av_readdata_pre[22] (
	.clk(clk),
	.d(\av_readdata_pre[22]~19_combout ),
	.asdata(b_full),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_22),
	.prn(vcc));
defparam \av_readdata_pre[22] .is_wysiwyg = "true";
defparam \av_readdata_pre[22] .power_up = "low";

dffeas \av_readdata_pre[21] (
	.clk(clk),
	.d(\av_readdata_pre[21]~17_combout ),
	.asdata(counter_reg_bit_5),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_21),
	.prn(vcc));
defparam \av_readdata_pre[21] .is_wysiwyg = "true";
defparam \av_readdata_pre[21] .power_up = "low";

cycloneive_lcell_comb \read_latency_shift_reg~0 (
	.dataa(rst1),
	.datab(d_read),
	.datac(gnd),
	.datad(read_accepted),
	.cin(gnd),
	.combout(read_latency_shift_reg),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hEEFF;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cycloneive_lcell_comb \read_latency_shift_reg~1 (
	.dataa(rst1),
	.datab(d_read),
	.datac(av_waitrequest),
	.datad(read_accepted),
	.cin(gnd),
	.combout(read_latency_shift_reg1),
	.cout());
defparam \read_latency_shift_reg~1 .lut_mask = 16'hFEFF;
defparam \read_latency_shift_reg~1 .sum_lutc_input = "datac";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[12] (
	.clk(clk),
	.d(av_readdata[12]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_12),
	.prn(vcc));
defparam \av_readdata_pre[12] .is_wysiwyg = "true";
defparam \av_readdata_pre[12] .power_up = "low";

dffeas \av_readdata_pre[10] (
	.clk(clk),
	.d(av_readdata[10]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_10),
	.prn(vcc));
defparam \av_readdata_pre[10] .is_wysiwyg = "true";
defparam \av_readdata_pre[10] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[15] (
	.clk(clk),
	.d(av_readdata[15]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_15),
	.prn(vcc));
defparam \av_readdata_pre[15] .is_wysiwyg = "true";
defparam \av_readdata_pre[15] .power_up = "low";

dffeas \av_readdata_pre[14] (
	.clk(clk),
	.d(av_readdata[14]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_14),
	.prn(vcc));
defparam \av_readdata_pre[14] .is_wysiwyg = "true";
defparam \av_readdata_pre[14] .power_up = "low";

dffeas \av_readdata_pre[13] (
	.clk(clk),
	.d(\av_readdata_pre[13]~21_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_13),
	.prn(vcc));
defparam \av_readdata_pre[13] .is_wysiwyg = "true";
defparam \av_readdata_pre[13] .power_up = "low";

cycloneive_lcell_comb \av_readdata_pre[16]~7 (
	.dataa(counter_reg_bit_01),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\av_readdata_pre[16]~7_combout ),
	.cout(\av_readdata_pre[16]~8 ));
defparam \av_readdata_pre[16]~7 .lut_mask = 16'hAA55;
defparam \av_readdata_pre[16]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata_pre[17]~9 (
	.dataa(counter_reg_bit_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\av_readdata_pre[16]~8 ),
	.combout(\av_readdata_pre[17]~9_combout ),
	.cout(\av_readdata_pre[17]~10 ));
defparam \av_readdata_pre[17]~9 .lut_mask = 16'h5AAF;
defparam \av_readdata_pre[17]~9 .sum_lutc_input = "cin";

cycloneive_lcell_comb \av_readdata_pre[18]~11 (
	.dataa(counter_reg_bit_21),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\av_readdata_pre[17]~10 ),
	.combout(\av_readdata_pre[18]~11_combout ),
	.cout(\av_readdata_pre[18]~12 ));
defparam \av_readdata_pre[18]~11 .lut_mask = 16'h5A5F;
defparam \av_readdata_pre[18]~11 .sum_lutc_input = "cin";

cycloneive_lcell_comb \av_readdata_pre[19]~13 (
	.dataa(counter_reg_bit_31),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\av_readdata_pre[18]~12 ),
	.combout(\av_readdata_pre[19]~13_combout ),
	.cout(\av_readdata_pre[19]~14 ));
defparam \av_readdata_pre[19]~13 .lut_mask = 16'h5AAF;
defparam \av_readdata_pre[19]~13 .sum_lutc_input = "cin";

cycloneive_lcell_comb \av_readdata_pre[20]~15 (
	.dataa(counter_reg_bit_41),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\av_readdata_pre[19]~14 ),
	.combout(\av_readdata_pre[20]~15_combout ),
	.cout(\av_readdata_pre[20]~16 ));
defparam \av_readdata_pre[20]~15 .lut_mask = 16'h5A5F;
defparam \av_readdata_pre[20]~15 .sum_lutc_input = "cin";

cycloneive_lcell_comb \av_readdata_pre[21]~17 (
	.dataa(counter_reg_bit_51),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\av_readdata_pre[20]~16 ),
	.combout(\av_readdata_pre[21]~17_combout ),
	.cout(\av_readdata_pre[21]~18 ));
defparam \av_readdata_pre[21]~17 .lut_mask = 16'h5AAF;
defparam \av_readdata_pre[21]~17 .sum_lutc_input = "cin";

cycloneive_lcell_comb \av_readdata_pre[22]~19 (
	.dataa(b_full1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\av_readdata_pre[21]~18 ),
	.combout(\av_readdata_pre[22]~19_combout ),
	.cout());
defparam \av_readdata_pre[22]~19 .lut_mask = 16'h5A5A;
defparam \av_readdata_pre[22]~19 .sum_lutc_input = "cin";

cycloneive_lcell_comb \read_latency_shift_reg~2 (
	.dataa(Equal3),
	.datab(read_latency_shift_reg1),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\read_latency_shift_reg~2_combout ),
	.cout());
defparam \read_latency_shift_reg~2 .lut_mask = 16'hEEFF;
defparam \read_latency_shift_reg~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_readdata_pre[13]~21 (
	.dataa(b_full1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\av_readdata_pre[13]~21_combout ),
	.cout());
defparam \av_readdata_pre[13]~21 .lut_mask = 16'h5555;
defparam \av_readdata_pre[13]~21 .sum_lutc_input = "datac";

endmodule

module nios_mcu_altera_merlin_slave_translator_2 (
	av_readdata,
	reset,
	rst1,
	read_latency_shift_reg_0,
	write,
	mem,
	WideOr1,
	av_readdata_pre_0,
	av_readdata_pre_22,
	av_readdata_pre_23,
	av_readdata_pre_24,
	av_readdata_pre_25,
	av_readdata_pre_26,
	av_readdata_pre_11,
	av_readdata_pre_13,
	av_readdata_pre_16,
	av_readdata_pre_12,
	av_readdata_pre_1,
	av_readdata_pre_3,
	av_readdata_pre_2,
	av_readdata_pre_5,
	av_readdata_pre_4,
	av_readdata_pre_14,
	av_readdata_pre_15,
	av_readdata_pre_18,
	av_readdata_pre_17,
	av_readdata_pre_10,
	av_readdata_pre_9,
	av_readdata_pre_8,
	av_readdata_pre_7,
	av_readdata_pre_6,
	av_readdata_pre_21,
	av_readdata_pre_19,
	av_readdata_pre_20,
	av_readdata_pre_27,
	av_readdata_pre_28,
	av_readdata_pre_29,
	av_readdata_pre_30,
	av_readdata_pre_31,
	clk)/* synthesis synthesis_greybox=1 */;
input 	[31:0] av_readdata;
input 	reset;
input 	rst1;
output 	read_latency_shift_reg_0;
input 	write;
input 	mem;
input 	WideOr1;
output 	av_readdata_pre_0;
output 	av_readdata_pre_22;
output 	av_readdata_pre_23;
output 	av_readdata_pre_24;
output 	av_readdata_pre_25;
output 	av_readdata_pre_26;
output 	av_readdata_pre_11;
output 	av_readdata_pre_13;
output 	av_readdata_pre_16;
output 	av_readdata_pre_12;
output 	av_readdata_pre_1;
output 	av_readdata_pre_3;
output 	av_readdata_pre_2;
output 	av_readdata_pre_5;
output 	av_readdata_pre_4;
output 	av_readdata_pre_14;
output 	av_readdata_pre_15;
output 	av_readdata_pre_18;
output 	av_readdata_pre_17;
output 	av_readdata_pre_10;
output 	av_readdata_pre_9;
output 	av_readdata_pre_8;
output 	av_readdata_pre_7;
output 	av_readdata_pre_6;
output 	av_readdata_pre_21;
output 	av_readdata_pre_19;
output 	av_readdata_pre_20;
output 	av_readdata_pre_27;
output 	av_readdata_pre_28;
output 	av_readdata_pre_29;
output 	av_readdata_pre_30;
output 	av_readdata_pre_31;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~0_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[22] (
	.clk(clk),
	.d(av_readdata[22]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_22),
	.prn(vcc));
defparam \av_readdata_pre[22] .is_wysiwyg = "true";
defparam \av_readdata_pre[22] .power_up = "low";

dffeas \av_readdata_pre[23] (
	.clk(clk),
	.d(av_readdata[23]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_23),
	.prn(vcc));
defparam \av_readdata_pre[23] .is_wysiwyg = "true";
defparam \av_readdata_pre[23] .power_up = "low";

dffeas \av_readdata_pre[24] (
	.clk(clk),
	.d(av_readdata[24]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_24),
	.prn(vcc));
defparam \av_readdata_pre[24] .is_wysiwyg = "true";
defparam \av_readdata_pre[24] .power_up = "low";

dffeas \av_readdata_pre[25] (
	.clk(clk),
	.d(av_readdata[25]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_25),
	.prn(vcc));
defparam \av_readdata_pre[25] .is_wysiwyg = "true";
defparam \av_readdata_pre[25] .power_up = "low";

dffeas \av_readdata_pre[26] (
	.clk(clk),
	.d(av_readdata[26]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_26),
	.prn(vcc));
defparam \av_readdata_pre[26] .is_wysiwyg = "true";
defparam \av_readdata_pre[26] .power_up = "low";

dffeas \av_readdata_pre[11] (
	.clk(clk),
	.d(av_readdata[11]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_11),
	.prn(vcc));
defparam \av_readdata_pre[11] .is_wysiwyg = "true";
defparam \av_readdata_pre[11] .power_up = "low";

dffeas \av_readdata_pre[13] (
	.clk(clk),
	.d(av_readdata[13]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_13),
	.prn(vcc));
defparam \av_readdata_pre[13] .is_wysiwyg = "true";
defparam \av_readdata_pre[13] .power_up = "low";

dffeas \av_readdata_pre[16] (
	.clk(clk),
	.d(av_readdata[16]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_16),
	.prn(vcc));
defparam \av_readdata_pre[16] .is_wysiwyg = "true";
defparam \av_readdata_pre[16] .power_up = "low";

dffeas \av_readdata_pre[12] (
	.clk(clk),
	.d(av_readdata[12]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_12),
	.prn(vcc));
defparam \av_readdata_pre[12] .is_wysiwyg = "true";
defparam \av_readdata_pre[12] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[14] (
	.clk(clk),
	.d(av_readdata[14]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_14),
	.prn(vcc));
defparam \av_readdata_pre[14] .is_wysiwyg = "true";
defparam \av_readdata_pre[14] .power_up = "low";

dffeas \av_readdata_pre[15] (
	.clk(clk),
	.d(av_readdata[15]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_15),
	.prn(vcc));
defparam \av_readdata_pre[15] .is_wysiwyg = "true";
defparam \av_readdata_pre[15] .power_up = "low";

dffeas \av_readdata_pre[18] (
	.clk(clk),
	.d(av_readdata[18]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_18),
	.prn(vcc));
defparam \av_readdata_pre[18] .is_wysiwyg = "true";
defparam \av_readdata_pre[18] .power_up = "low";

dffeas \av_readdata_pre[17] (
	.clk(clk),
	.d(av_readdata[17]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_17),
	.prn(vcc));
defparam \av_readdata_pre[17] .is_wysiwyg = "true";
defparam \av_readdata_pre[17] .power_up = "low";

dffeas \av_readdata_pre[10] (
	.clk(clk),
	.d(av_readdata[10]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_10),
	.prn(vcc));
defparam \av_readdata_pre[10] .is_wysiwyg = "true";
defparam \av_readdata_pre[10] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[21] (
	.clk(clk),
	.d(av_readdata[21]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_21),
	.prn(vcc));
defparam \av_readdata_pre[21] .is_wysiwyg = "true";
defparam \av_readdata_pre[21] .power_up = "low";

dffeas \av_readdata_pre[19] (
	.clk(clk),
	.d(av_readdata[19]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_19),
	.prn(vcc));
defparam \av_readdata_pre[19] .is_wysiwyg = "true";
defparam \av_readdata_pre[19] .power_up = "low";

dffeas \av_readdata_pre[20] (
	.clk(clk),
	.d(av_readdata[20]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_20),
	.prn(vcc));
defparam \av_readdata_pre[20] .is_wysiwyg = "true";
defparam \av_readdata_pre[20] .power_up = "low";

dffeas \av_readdata_pre[27] (
	.clk(clk),
	.d(av_readdata[27]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_27),
	.prn(vcc));
defparam \av_readdata_pre[27] .is_wysiwyg = "true";
defparam \av_readdata_pre[27] .power_up = "low";

dffeas \av_readdata_pre[28] (
	.clk(clk),
	.d(av_readdata[28]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_28),
	.prn(vcc));
defparam \av_readdata_pre[28] .is_wysiwyg = "true";
defparam \av_readdata_pre[28] .power_up = "low";

dffeas \av_readdata_pre[29] (
	.clk(clk),
	.d(av_readdata[29]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_29),
	.prn(vcc));
defparam \av_readdata_pre[29] .is_wysiwyg = "true";
defparam \av_readdata_pre[29] .power_up = "low";

dffeas \av_readdata_pre[30] (
	.clk(clk),
	.d(av_readdata[30]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_30),
	.prn(vcc));
defparam \av_readdata_pre[30] .is_wysiwyg = "true";
defparam \av_readdata_pre[30] .power_up = "low";

dffeas \av_readdata_pre[31] (
	.clk(clk),
	.d(av_readdata[31]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_31),
	.prn(vcc));
defparam \av_readdata_pre[31] .is_wysiwyg = "true";
defparam \av_readdata_pre[31] .power_up = "low";

cycloneive_lcell_comb \read_latency_shift_reg~0 (
	.dataa(rst1),
	.datab(write),
	.datac(WideOr1),
	.datad(mem),
	.cin(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hFFFE;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

endmodule

module nios_mcu_altera_merlin_slave_translator_3 (
	reset,
	rst1,
	F_pc_9,
	read_accepted,
	i_read,
	read_latency_shift_reg,
	Equal0,
	read_latency_shift_reg_0,
	mem_used_1,
	read_latency_shift_reg1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	rst1;
input 	F_pc_9;
input 	read_accepted;
input 	i_read;
output 	read_latency_shift_reg;
input 	Equal0;
output 	read_latency_shift_reg_0;
input 	mem_used_1;
output 	read_latency_shift_reg1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \read_latency_shift_reg~0 (
	.dataa(rst1),
	.datab(gnd),
	.datac(read_accepted),
	.datad(i_read),
	.cin(gnd),
	.combout(read_latency_shift_reg),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hAFFF;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(read_latency_shift_reg1),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cycloneive_lcell_comb \read_latency_shift_reg~1 (
	.dataa(read_latency_shift_reg),
	.datab(F_pc_9),
	.datac(Equal0),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(read_latency_shift_reg1),
	.cout());
defparam \read_latency_shift_reg~1 .lut_mask = 16'hBFFF;
defparam \read_latency_shift_reg~1 .sum_lutc_input = "datac";

endmodule

module nios_mcu_altera_merlin_slave_translator_4 (
	reset,
	read_latency_shift_reg,
	read_latency_shift_reg_0,
	src_channel_4,
	mem_used_1,
	read_latency_shift_reg1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	read_latency_shift_reg;
output 	read_latency_shift_reg_0;
input 	src_channel_4;
input 	mem_used_1;
output 	read_latency_shift_reg1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(read_latency_shift_reg1),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cycloneive_lcell_comb \read_latency_shift_reg~0 (
	.dataa(read_latency_shift_reg),
	.datab(src_channel_4),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(read_latency_shift_reg1),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hEEFF;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

endmodule

module nios_mcu_altera_merlin_slave_translator_5 (
	W_alu_result_4,
	reset,
	Equal1,
	mem_used_1,
	always0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	read_latency_shift_reg_0,
	read_latency_shift_reg,
	Equal11,
	m0_write,
	wait_latency_counter_11,
	read_latency_shift_reg1,
	always2,
	read_latency_shift_reg2,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata,
	clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_4;
input 	reset;
input 	Equal1;
input 	mem_used_1;
input 	always0;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
output 	read_latency_shift_reg_0;
input 	read_latency_shift_reg;
input 	Equal11;
input 	m0_write;
output 	wait_latency_counter_11;
output 	read_latency_shift_reg1;
input 	always2;
output 	read_latency_shift_reg2;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~0_combout ;
wire \wait_latency_counter~1_combout ;
wire \wait_latency_counter~2_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(read_latency_shift_reg2),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cycloneive_lcell_comb \wait_latency_counter[1]~0 (
	.dataa(wait_latency_counter_0),
	.datab(always0),
	.datac(m0_write),
	.datad(wait_latency_counter_1),
	.cin(gnd),
	.combout(wait_latency_counter_11),
	.cout());
defparam \wait_latency_counter[1]~0 .lut_mask = 16'h96FF;
defparam \wait_latency_counter[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_latency_shift_reg~0 (
	.dataa(Equal1),
	.datab(wait_latency_counter_11),
	.datac(W_alu_result_4),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(read_latency_shift_reg1),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hEFFF;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_latency_shift_reg~1 (
	.dataa(Equal11),
	.datab(wait_latency_counter_11),
	.datac(read_latency_shift_reg),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(read_latency_shift_reg2),
	.cout());
defparam \read_latency_shift_reg~1 .lut_mask = 16'hFEFF;
defparam \read_latency_shift_reg~1 .sum_lutc_input = "datac";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

cycloneive_lcell_comb \Add0~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(wait_latency_counter_1),
	.datad(wait_latency_counter_0),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout());
defparam \Add0~0 .lut_mask = 16'h0FF0;
defparam \Add0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wait_latency_counter~1 (
	.dataa(always0),
	.datab(always2),
	.datac(\Add0~0_combout ),
	.datad(wait_latency_counter_11),
	.cin(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.cout());
defparam \wait_latency_counter~1 .lut_mask = 16'hFEFF;
defparam \wait_latency_counter~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wait_latency_counter~2 (
	.dataa(wait_latency_counter_0),
	.datab(wait_latency_counter_11),
	.datac(always0),
	.datad(always2),
	.cin(gnd),
	.combout(\wait_latency_counter~2_combout ),
	.cout());
defparam \wait_latency_counter~2 .lut_mask = 16'hFFF7;
defparam \wait_latency_counter~2 .sum_lutc_input = "datac";

endmodule

module nios_mcu_nios_mcu_mm_interconnect_0_cmd_demux (
	W_alu_result_11,
	rst1,
	Equal0,
	Equal3,
	src_channel_4,
	mem_used_1,
	sink_ready,
	saved_grant_0,
	write,
	av_waitrequest,
	mem_used_11,
	WideOr0,
	Equal2,
	dRead,
	always2,
	mem_used_12,
	sReadCountPipelined_0,
	sink_ready1,
	WideOr01,
	src2_valid)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_11;
input 	rst1;
input 	Equal0;
input 	Equal3;
input 	src_channel_4;
input 	mem_used_1;
output 	sink_ready;
input 	saved_grant_0;
input 	write;
input 	av_waitrequest;
input 	mem_used_11;
output 	WideOr0;
input 	Equal2;
input 	dRead;
input 	always2;
input 	mem_used_12;
input 	sReadCountPipelined_0;
output 	sink_ready1;
output 	WideOr01;
output 	src2_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \sink_ready~1_combout ;


cycloneive_lcell_comb \sink_ready~0 (
	.dataa(rst1),
	.datab(src_channel_4),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(sink_ready),
	.cout());
defparam \sink_ready~0 .lut_mask = 16'hEEFF;
defparam \sink_ready~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~0 (
	.dataa(\sink_ready~1_combout ),
	.datab(Equal3),
	.datac(av_waitrequest),
	.datad(mem_used_11),
	.cin(gnd),
	.combout(WideOr0),
	.cout());
defparam \WideOr0~0 .lut_mask = 16'hFEFF;
defparam \WideOr0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sink_ready~2 (
	.dataa(Equal2),
	.datab(dRead),
	.datac(sReadCountPipelined_0),
	.datad(mem_used_12),
	.cin(gnd),
	.combout(sink_ready1),
	.cout());
defparam \sink_ready~2 .lut_mask = 16'hEFFF;
defparam \sink_ready~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~1 (
	.dataa(WideOr0),
	.datab(rst1),
	.datac(src_channel_4),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(WideOr01),
	.cout());
defparam \WideOr0~1 .lut_mask = 16'hFEFF;
defparam \WideOr0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src2_valid~0 (
	.dataa(W_alu_result_11),
	.datab(rst1),
	.datac(always2),
	.datad(Equal0),
	.cin(gnd),
	.combout(src2_valid),
	.cout());
defparam \src2_valid~0 .lut_mask = 16'hFEFF;
defparam \src2_valid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sink_ready~1 (
	.dataa(W_alu_result_11),
	.datab(saved_grant_0),
	.datac(write),
	.datad(Equal0),
	.cin(gnd),
	.combout(\sink_ready~1_combout ),
	.cout());
defparam \sink_ready~1 .lut_mask = 16'hFEFF;
defparam \sink_ready~1 .sum_lutc_input = "datac";

endmodule

module nios_mcu_nios_mcu_mm_interconnect_0_cmd_demux_001 (
	F_pc_9,
	read_latency_shift_reg,
	Equal0,
	src0_valid)/* synthesis synthesis_greybox=1 */;
input 	F_pc_9;
input 	read_latency_shift_reg;
input 	Equal0;
output 	src0_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \src0_valid~0 (
	.dataa(F_pc_9),
	.datab(read_latency_shift_reg),
	.datac(Equal0),
	.datad(gnd),
	.cin(gnd),
	.combout(src0_valid),
	.cout());
defparam \src0_valid~0 .lut_mask = 16'hFEFE;
defparam \src0_valid~0 .sum_lutc_input = "datac";

endmodule

module nios_mcu_nios_mcu_mm_interconnect_0_cmd_demux_001_1 (
	mem_73_0,
	mem_55_0,
	read_latency_shift_reg_0,
	src0_valid,
	src1_valid)/* synthesis synthesis_greybox=1 */;
input 	mem_73_0;
input 	mem_55_0;
input 	read_latency_shift_reg_0;
output 	src0_valid;
output 	src1_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \src0_valid~0 (
	.dataa(read_latency_shift_reg_0),
	.datab(gnd),
	.datac(mem_73_0),
	.datad(mem_55_0),
	.cin(gnd),
	.combout(src0_valid),
	.cout());
defparam \src0_valid~0 .lut_mask = 16'hAFFF;
defparam \src0_valid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src1_valid~0 (
	.dataa(read_latency_shift_reg_0),
	.datab(mem_73_0),
	.datac(mem_55_0),
	.datad(gnd),
	.cin(gnd),
	.combout(src1_valid),
	.cout());
defparam \src1_valid~0 .lut_mask = 16'hFEFE;
defparam \src1_valid~0 .sum_lutc_input = "datac";

endmodule

module nios_mcu_nios_mcu_mm_interconnect_0_cmd_mux_002 (
	W_alu_result_10,
	W_alu_result_9,
	W_alu_result_8,
	W_alu_result_7,
	W_alu_result_6,
	W_alu_result_5,
	W_alu_result_4,
	W_alu_result_3,
	W_alu_result_2,
	d_writedata_24,
	d_writedata_25,
	d_writedata_26,
	d_writedata_27,
	d_writedata_28,
	d_writedata_29,
	d_writedata_30,
	d_writedata_31,
	d_writedata_0,
	r_sync_rst,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	saved_grant_0,
	waitrequest,
	mem_used_1,
	F_pc_8,
	F_pc_7,
	F_pc_6,
	F_pc_5,
	F_pc_4,
	F_pc_3,
	F_pc_2,
	F_pc_1,
	F_pc_0,
	saved_grant_1,
	src0_valid,
	src2_valid,
	WideOr11,
	hbreak_enabled,
	src_data_46,
	d_byteenable_0,
	d_writedata_22,
	d_byteenable_2,
	d_writedata_23,
	d_byteenable_3,
	d_writedata_11,
	d_byteenable_1,
	d_writedata_13,
	d_writedata_16,
	d_writedata_12,
	d_writedata_14,
	d_writedata_15,
	d_writedata_18,
	d_writedata_17,
	d_writedata_10,
	d_writedata_9,
	d_writedata_8,
	d_writedata_21,
	d_writedata_19,
	d_writedata_20,
	src_payload,
	src_payload1,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_32,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_data_34,
	src_payload6,
	src_payload7,
	src_data_35,
	src_payload8,
	src_payload9,
	src_payload10,
	src_data_33,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_10;
input 	W_alu_result_9;
input 	W_alu_result_8;
input 	W_alu_result_7;
input 	W_alu_result_6;
input 	W_alu_result_5;
input 	W_alu_result_4;
input 	W_alu_result_3;
input 	W_alu_result_2;
input 	d_writedata_24;
input 	d_writedata_25;
input 	d_writedata_26;
input 	d_writedata_27;
input 	d_writedata_28;
input 	d_writedata_29;
input 	d_writedata_30;
input 	d_writedata_31;
input 	d_writedata_0;
input 	r_sync_rst;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	d_writedata_6;
input 	d_writedata_7;
output 	saved_grant_0;
input 	waitrequest;
input 	mem_used_1;
input 	F_pc_8;
input 	F_pc_7;
input 	F_pc_6;
input 	F_pc_5;
input 	F_pc_4;
input 	F_pc_3;
input 	F_pc_2;
input 	F_pc_1;
input 	F_pc_0;
output 	saved_grant_1;
input 	src0_valid;
input 	src2_valid;
output 	WideOr11;
input 	hbreak_enabled;
output 	src_data_46;
input 	d_byteenable_0;
input 	d_writedata_22;
input 	d_byteenable_2;
input 	d_writedata_23;
input 	d_byteenable_3;
input 	d_writedata_11;
input 	d_byteenable_1;
input 	d_writedata_13;
input 	d_writedata_16;
input 	d_writedata_12;
input 	d_writedata_14;
input 	d_writedata_15;
input 	d_writedata_18;
input 	d_writedata_17;
input 	d_writedata_10;
input 	d_writedata_9;
input 	d_writedata_8;
input 	d_writedata_21;
input 	d_writedata_19;
input 	d_writedata_20;
output 	src_payload;
output 	src_payload1;
output 	src_data_38;
output 	src_data_39;
output 	src_data_40;
output 	src_data_41;
output 	src_data_42;
output 	src_data_43;
output 	src_data_44;
output 	src_data_45;
output 	src_data_32;
output 	src_payload2;
output 	src_payload3;
output 	src_payload4;
output 	src_payload5;
output 	src_data_34;
output 	src_payload6;
output 	src_payload7;
output 	src_data_35;
output 	src_payload8;
output 	src_payload9;
output 	src_payload10;
output 	src_data_33;
output 	src_payload11;
output 	src_payload12;
output 	src_payload13;
output 	src_payload14;
output 	src_payload15;
output 	src_payload16;
output 	src_payload17;
output 	src_payload18;
output 	src_payload19;
output 	src_payload20;
output 	src_payload21;
output 	src_payload22;
output 	src_payload23;
output 	src_payload24;
output 	src_payload25;
output 	src_payload26;
output 	src_payload27;
output 	src_payload28;
output 	src_payload29;
output 	src_payload30;
output 	src_payload31;
output 	src_payload32;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[0]~0_combout ;
wire \arb|grant[1]~1_combout ;
wire \update_grant~0_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~1_combout ;


nios_mcu_altera_merlin_arbitrator arb(
	.reset(r_sync_rst),
	.src0_valid(src0_valid),
	.src2_valid(src2_valid),
	.grant_0(\arb|grant[0]~0_combout ),
	.update_grant(\update_grant~1_combout ),
	.grant_1(\arb|grant[1]~1_combout ),
	.clk(clk_clk));

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~1_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~1_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cycloneive_lcell_comb WideOr1(
	.dataa(saved_grant_0),
	.datab(src0_valid),
	.datac(saved_grant_1),
	.datad(src2_valid),
	.cin(gnd),
	.combout(WideOr11),
	.cout());
defparam WideOr1.lut_mask = 16'hFFFE;
defparam WideOr1.sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[46] (
	.dataa(W_alu_result_10),
	.datab(F_pc_8),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_46),
	.cout());
defparam \src_data[46] .lut_mask = 16'hFFFE;
defparam \src_data[46] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~0 (
	.dataa(saved_grant_0),
	.datab(hbreak_enabled),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload),
	.cout());
defparam \src_payload~0 .lut_mask = 16'hEEEE;
defparam \src_payload~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~1 (
	.dataa(d_writedata_0),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload1),
	.cout());
defparam \src_payload~1 .lut_mask = 16'hEEEE;
defparam \src_payload~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[38] (
	.dataa(W_alu_result_2),
	.datab(F_pc_0),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_38),
	.cout());
defparam \src_data[38] .lut_mask = 16'hFFFE;
defparam \src_data[38] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[39] (
	.dataa(W_alu_result_3),
	.datab(F_pc_1),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_39),
	.cout());
defparam \src_data[39] .lut_mask = 16'hFFFE;
defparam \src_data[39] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[40] (
	.dataa(W_alu_result_4),
	.datab(F_pc_2),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_40),
	.cout());
defparam \src_data[40] .lut_mask = 16'hFFFE;
defparam \src_data[40] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[41] (
	.dataa(W_alu_result_5),
	.datab(F_pc_3),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_41),
	.cout());
defparam \src_data[41] .lut_mask = 16'hFFFE;
defparam \src_data[41] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[42] (
	.dataa(W_alu_result_6),
	.datab(F_pc_4),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_42),
	.cout());
defparam \src_data[42] .lut_mask = 16'hFFFE;
defparam \src_data[42] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[43] (
	.dataa(W_alu_result_7),
	.datab(F_pc_5),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_43),
	.cout());
defparam \src_data[43] .lut_mask = 16'hFFFE;
defparam \src_data[43] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[44] (
	.dataa(W_alu_result_8),
	.datab(F_pc_6),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_44),
	.cout());
defparam \src_data[44] .lut_mask = 16'hFFFE;
defparam \src_data[44] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[45] (
	.dataa(W_alu_result_9),
	.datab(F_pc_7),
	.datac(saved_grant_1),
	.datad(saved_grant_0),
	.cin(gnd),
	.combout(src_data_45),
	.cout());
defparam \src_data[45] .lut_mask = 16'hFFFE;
defparam \src_data[45] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[32] (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(d_byteenable_0),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_32),
	.cout());
defparam \src_data[32] .lut_mask = 16'hFEFE;
defparam \src_data[32] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~2 (
	.dataa(d_writedata_1),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload2),
	.cout());
defparam \src_payload~2 .lut_mask = 16'hEEEE;
defparam \src_payload~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~3 (
	.dataa(d_writedata_3),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload3),
	.cout());
defparam \src_payload~3 .lut_mask = 16'hEEEE;
defparam \src_payload~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~4 (
	.dataa(d_writedata_2),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload4),
	.cout());
defparam \src_payload~4 .lut_mask = 16'hEEEE;
defparam \src_payload~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~5 (
	.dataa(saved_grant_0),
	.datab(d_writedata_22),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload5),
	.cout());
defparam \src_payload~5 .lut_mask = 16'hEEEE;
defparam \src_payload~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[34] (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(d_byteenable_2),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_34),
	.cout());
defparam \src_data[34] .lut_mask = 16'hFEFE;
defparam \src_data[34] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~6 (
	.dataa(saved_grant_0),
	.datab(d_writedata_23),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload6),
	.cout());
defparam \src_payload~6 .lut_mask = 16'hEEEE;
defparam \src_payload~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~7 (
	.dataa(saved_grant_0),
	.datab(d_writedata_24),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload7),
	.cout());
defparam \src_payload~7 .lut_mask = 16'hEEEE;
defparam \src_payload~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[35] (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(d_byteenable_3),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_35),
	.cout());
defparam \src_data[35] .lut_mask = 16'hFEFE;
defparam \src_data[35] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~8 (
	.dataa(saved_grant_0),
	.datab(d_writedata_25),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload8),
	.cout());
defparam \src_payload~8 .lut_mask = 16'hEEEE;
defparam \src_payload~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~9 (
	.dataa(saved_grant_0),
	.datab(d_writedata_26),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload9),
	.cout());
defparam \src_payload~9 .lut_mask = 16'hEEEE;
defparam \src_payload~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~10 (
	.dataa(saved_grant_0),
	.datab(d_writedata_11),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload10),
	.cout());
defparam \src_payload~10 .lut_mask = 16'hEEEE;
defparam \src_payload~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[33] (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(d_byteenable_1),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_33),
	.cout());
defparam \src_data[33] .lut_mask = 16'hFEFE;
defparam \src_data[33] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~11 (
	.dataa(saved_grant_0),
	.datab(d_writedata_13),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload11),
	.cout());
defparam \src_payload~11 .lut_mask = 16'hEEEE;
defparam \src_payload~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~12 (
	.dataa(saved_grant_0),
	.datab(d_writedata_16),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload12),
	.cout());
defparam \src_payload~12 .lut_mask = 16'hEEEE;
defparam \src_payload~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~13 (
	.dataa(saved_grant_0),
	.datab(d_writedata_12),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload13),
	.cout());
defparam \src_payload~13 .lut_mask = 16'hEEEE;
defparam \src_payload~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~14 (
	.dataa(d_writedata_5),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload14),
	.cout());
defparam \src_payload~14 .lut_mask = 16'hEEEE;
defparam \src_payload~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~15 (
	.dataa(d_writedata_4),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload15),
	.cout());
defparam \src_payload~15 .lut_mask = 16'hEEEE;
defparam \src_payload~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~16 (
	.dataa(saved_grant_0),
	.datab(d_writedata_14),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload16),
	.cout());
defparam \src_payload~16 .lut_mask = 16'hEEEE;
defparam \src_payload~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~17 (
	.dataa(saved_grant_0),
	.datab(d_writedata_15),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload17),
	.cout());
defparam \src_payload~17 .lut_mask = 16'hEEEE;
defparam \src_payload~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~18 (
	.dataa(saved_grant_0),
	.datab(d_writedata_18),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload18),
	.cout());
defparam \src_payload~18 .lut_mask = 16'hEEEE;
defparam \src_payload~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~19 (
	.dataa(saved_grant_0),
	.datab(d_writedata_17),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload19),
	.cout());
defparam \src_payload~19 .lut_mask = 16'hEEEE;
defparam \src_payload~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~20 (
	.dataa(saved_grant_0),
	.datab(d_writedata_10),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload20),
	.cout());
defparam \src_payload~20 .lut_mask = 16'hEEEE;
defparam \src_payload~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~21 (
	.dataa(saved_grant_0),
	.datab(d_writedata_9),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload21),
	.cout());
defparam \src_payload~21 .lut_mask = 16'hEEEE;
defparam \src_payload~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~22 (
	.dataa(saved_grant_0),
	.datab(d_writedata_8),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload22),
	.cout());
defparam \src_payload~22 .lut_mask = 16'hEEEE;
defparam \src_payload~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~23 (
	.dataa(d_writedata_7),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload23),
	.cout());
defparam \src_payload~23 .lut_mask = 16'hEEEE;
defparam \src_payload~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~24 (
	.dataa(d_writedata_6),
	.datab(saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload24),
	.cout());
defparam \src_payload~24 .lut_mask = 16'hEEEE;
defparam \src_payload~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~25 (
	.dataa(saved_grant_0),
	.datab(d_writedata_21),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload25),
	.cout());
defparam \src_payload~25 .lut_mask = 16'hEEEE;
defparam \src_payload~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~26 (
	.dataa(saved_grant_0),
	.datab(d_writedata_19),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload26),
	.cout());
defparam \src_payload~26 .lut_mask = 16'hEEEE;
defparam \src_payload~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~27 (
	.dataa(saved_grant_0),
	.datab(d_writedata_20),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload27),
	.cout());
defparam \src_payload~27 .lut_mask = 16'hEEEE;
defparam \src_payload~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~28 (
	.dataa(saved_grant_0),
	.datab(d_writedata_27),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload28),
	.cout());
defparam \src_payload~28 .lut_mask = 16'hEEEE;
defparam \src_payload~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~29 (
	.dataa(saved_grant_0),
	.datab(d_writedata_28),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload29),
	.cout());
defparam \src_payload~29 .lut_mask = 16'hEEEE;
defparam \src_payload~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~30 (
	.dataa(saved_grant_0),
	.datab(d_writedata_29),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload30),
	.cout());
defparam \src_payload~30 .lut_mask = 16'hEEEE;
defparam \src_payload~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~31 (
	.dataa(saved_grant_0),
	.datab(d_writedata_30),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload31),
	.cout());
defparam \src_payload~31 .lut_mask = 16'hEEEE;
defparam \src_payload~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~32 (
	.dataa(saved_grant_0),
	.datab(d_writedata_31),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload32),
	.cout());
defparam \src_payload~32 .lut_mask = 16'hEEEE;
defparam \src_payload~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \update_grant~0 (
	.dataa(saved_grant_0),
	.datab(saved_grant_1),
	.datac(waitrequest),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\update_grant~0_combout ),
	.cout());
defparam \update_grant~0 .lut_mask = 16'hEFFF;
defparam \update_grant~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \packet_in_progress~0 (
	.dataa(\update_grant~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\packet_in_progress~0_combout ),
	.cout());
defparam \packet_in_progress~0 .lut_mask = 16'h5555;
defparam \packet_in_progress~0 .sum_lutc_input = "datac";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cycloneive_lcell_comb \update_grant~1 (
	.dataa(\update_grant~0_combout ),
	.datab(WideOr11),
	.datac(gnd),
	.datad(\packet_in_progress~q ),
	.cin(gnd),
	.combout(\update_grant~1_combout ),
	.cout());
defparam \update_grant~1 .lut_mask = 16'h88BB;
defparam \update_grant~1 .sum_lutc_input = "datac";

endmodule

module nios_mcu_altera_merlin_arbitrator (
	reset,
	src0_valid,
	src2_valid,
	grant_0,
	update_grant,
	grant_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	src0_valid;
input 	src2_valid;
output 	grant_0;
input 	update_grant;
output 	grant_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[0]~q ;


cycloneive_lcell_comb \grant[0]~0 (
	.dataa(src2_valid),
	.datab(\top_priority_reg[1]~q ),
	.datac(src0_valid),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_0),
	.cout());
defparam \grant[0]~0 .lut_mask = 16'hEFFF;
defparam \grant[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \grant[1]~1 (
	.dataa(src0_valid),
	.datab(\top_priority_reg[1]~q ),
	.datac(src2_valid),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_1),
	.cout());
defparam \grant[1]~1 .lut_mask = 16'hEFFF;
defparam \grant[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \top_priority_reg[0]~0 (
	.dataa(update_grant),
	.datab(src2_valid),
	.datac(src0_valid),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.cout());
defparam \top_priority_reg[0]~0 .lut_mask = 16'hFEFE;
defparam \top_priority_reg[0]~0 .sum_lutc_input = "datac";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cycloneive_lcell_comb \top_priority_reg[0]~1 (
	.dataa(grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.cout());
defparam \top_priority_reg[0]~1 .lut_mask = 16'h5555;
defparam \top_priority_reg[0]~1 .sum_lutc_input = "datac";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module nios_mcu_nios_mcu_mm_interconnect_0_router (
	W_alu_result_12,
	W_alu_result_15,
	W_alu_result_14,
	W_alu_result_13,
	W_alu_result_11,
	W_alu_result_10,
	W_alu_result_9,
	W_alu_result_8,
	W_alu_result_7,
	W_alu_result_6,
	W_alu_result_5,
	W_alu_result_4,
	W_alu_result_3,
	Equal1,
	Equal11,
	Equal0,
	Equal3,
	src_channel_4,
	Equal2)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_12;
input 	W_alu_result_15;
input 	W_alu_result_14;
input 	W_alu_result_13;
input 	W_alu_result_11;
input 	W_alu_result_10;
input 	W_alu_result_9;
input 	W_alu_result_8;
input 	W_alu_result_7;
input 	W_alu_result_6;
input 	W_alu_result_5;
input 	W_alu_result_4;
input 	W_alu_result_3;
output 	Equal1;
output 	Equal11;
output 	Equal0;
output 	Equal3;
output 	src_channel_4;
output 	Equal2;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Equal1~0_combout ;
wire \Equal1~1_combout ;
wire \Equal1~2_combout ;
wire \Equal3~0_combout ;


cycloneive_lcell_comb \Equal1~3 (
	.dataa(\Equal1~0_combout ),
	.datab(\Equal1~1_combout ),
	.datac(\Equal1~2_combout ),
	.datad(W_alu_result_5),
	.cin(gnd),
	.combout(Equal1),
	.cout());
defparam \Equal1~3 .lut_mask = 16'hFEFF;
defparam \Equal1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal1~4 (
	.dataa(Equal1),
	.datab(gnd),
	.datac(gnd),
	.datad(W_alu_result_4),
	.cin(gnd),
	.combout(Equal11),
	.cout());
defparam \Equal1~4 .lut_mask = 16'hAAFF;
defparam \Equal1~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~0 (
	.dataa(W_alu_result_12),
	.datab(W_alu_result_14),
	.datac(W_alu_result_13),
	.datad(W_alu_result_15),
	.cin(gnd),
	.combout(Equal0),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hFEFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal3~1 (
	.dataa(\Equal1~0_combout ),
	.datab(\Equal1~1_combout ),
	.datac(\Equal1~2_combout ),
	.datad(\Equal3~0_combout ),
	.cin(gnd),
	.combout(Equal3),
	.cout());
defparam \Equal3~1 .lut_mask = 16'hFFFE;
defparam \Equal3~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_channel[4]~0 (
	.dataa(Equal0),
	.datab(W_alu_result_11),
	.datac(Equal1),
	.datad(Equal3),
	.cin(gnd),
	.combout(src_channel_4),
	.cout());
defparam \src_channel[4]~0 .lut_mask = 16'hBFFF;
defparam \src_channel[4]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal2~0 (
	.dataa(W_alu_result_4),
	.datab(Equal1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(Equal2),
	.cout());
defparam \Equal2~0 .lut_mask = 16'hEEEE;
defparam \Equal2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal1~0 (
	.dataa(W_alu_result_12),
	.datab(W_alu_result_15),
	.datac(W_alu_result_14),
	.datad(W_alu_result_13),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
defparam \Equal1~0 .lut_mask = 16'hEFFF;
defparam \Equal1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal1~1 (
	.dataa(W_alu_result_11),
	.datab(W_alu_result_10),
	.datac(W_alu_result_9),
	.datad(W_alu_result_8),
	.cin(gnd),
	.combout(\Equal1~1_combout ),
	.cout());
defparam \Equal1~1 .lut_mask = 16'h7FFF;
defparam \Equal1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal1~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(W_alu_result_7),
	.datad(W_alu_result_6),
	.cin(gnd),
	.combout(\Equal1~2_combout ),
	.cout());
defparam \Equal1~2 .lut_mask = 16'h0FFF;
defparam \Equal1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal3~0 (
	.dataa(W_alu_result_5),
	.datab(gnd),
	.datac(W_alu_result_4),
	.datad(W_alu_result_3),
	.cin(gnd),
	.combout(\Equal3~0_combout ),
	.cout());
defparam \Equal3~0 .lut_mask = 16'hAFFF;
defparam \Equal3~0 .sum_lutc_input = "datac";

endmodule

module nios_mcu_nios_mcu_mm_interconnect_0_router_001 (
	F_pc_10,
	F_pc_9,
	F_pc_13,
	F_pc_12,
	F_pc_11,
	Equal0,
	Equal01)/* synthesis synthesis_greybox=1 */;
input 	F_pc_10;
input 	F_pc_9;
input 	F_pc_13;
input 	F_pc_12;
input 	F_pc_11;
output 	Equal0;
output 	Equal01;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \Equal0~0 (
	.dataa(F_pc_13),
	.datab(F_pc_10),
	.datac(F_pc_12),
	.datad(F_pc_11),
	.cin(gnd),
	.combout(Equal0),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hBFFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~1 (
	.dataa(F_pc_9),
	.datab(Equal0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(Equal01),
	.cout());
defparam \Equal0~1 .lut_mask = 16'hEEEE;
defparam \Equal0~1 .sum_lutc_input = "datac";

endmodule

module nios_mcu_nios_mcu_mm_interconnect_0_rsp_mux (
	q_b_22,
	q_b_23,
	q_b_11,
	q_b_13,
	q_b_16,
	q_b_12,
	q_b_14,
	q_b_15,
	q_b_18,
	q_b_17,
	q_b_10,
	q_b_9,
	q_b_8,
	q_b_21,
	q_b_19,
	q_b_20,
	av_readdata_pre_16,
	av_readdata_pre_20,
	av_readdata_pre_19,
	av_readdata_pre_18,
	av_readdata_pre_17,
	av_readdata_pre_22,
	av_readdata_pre_21,
	read_latency_shift_reg_0,
	mem_73_0,
	mem_55_0,
	read_latency_shift_reg_01,
	read_latency_shift_reg_02,
	WideOr11,
	read_latency_shift_reg_03,
	read_latency_shift_reg_04,
	WideOr12,
	WideOr13,
	src0_valid,
	av_readdata_pre_221,
	av_readdata_pre_23,
	av_readdata_pre_11,
	av_readdata_pre_13,
	av_readdata_pre_161,
	av_readdata_pre_12,
	av_readdata_pre_14,
	av_readdata_pre_15,
	av_readdata_pre_181,
	av_readdata_pre_171,
	av_readdata_pre_10,
	av_readdata_pre_9,
	av_readdata_pre_8,
	av_readdata_pre_211,
	av_readdata_pre_191,
	av_readdata_pre_201,
	av_readdata_pre_81,
	av_readdata_pre_82,
	src_data_8,
	av_readdata_pre_121,
	av_readdata_pre_122,
	src_data_12,
	av_readdata_pre_111,
	src_data_11,
	av_readdata_pre_101,
	av_readdata_pre_102,
	src_data_10,
	av_readdata_pre_91,
	av_readdata_pre_92,
	src_data_9,
	av_readdata_pre_151,
	av_readdata_pre_152,
	src_data_15,
	av_readdata_pre_141,
	av_readdata_pre_142,
	src_data_14,
	av_readdata_pre_131,
	av_readdata_pre_132,
	src_data_13,
	av_readdata_pre_162,
	src_data_16,
	av_readdata_pre_202,
	src_data_20,
	av_readdata_pre_192,
	src_data_19,
	av_readdata_pre_182,
	src_data_18,
	av_readdata_pre_172,
	src_data_17,
	av_readdata_pre_231,
	src_data_23,
	av_readdata_pre_222,
	src_data_22,
	av_readdata_pre_212,
	src_data_21)/* synthesis synthesis_greybox=1 */;
input 	q_b_22;
input 	q_b_23;
input 	q_b_11;
input 	q_b_13;
input 	q_b_16;
input 	q_b_12;
input 	q_b_14;
input 	q_b_15;
input 	q_b_18;
input 	q_b_17;
input 	q_b_10;
input 	q_b_9;
input 	q_b_8;
input 	q_b_21;
input 	q_b_19;
input 	q_b_20;
input 	av_readdata_pre_16;
input 	av_readdata_pre_20;
input 	av_readdata_pre_19;
input 	av_readdata_pre_18;
input 	av_readdata_pre_17;
input 	av_readdata_pre_22;
input 	av_readdata_pre_21;
input 	read_latency_shift_reg_0;
input 	mem_73_0;
input 	mem_55_0;
input 	read_latency_shift_reg_01;
input 	read_latency_shift_reg_02;
output 	WideOr11;
input 	read_latency_shift_reg_03;
input 	read_latency_shift_reg_04;
output 	WideOr12;
output 	WideOr13;
input 	src0_valid;
input 	av_readdata_pre_221;
input 	av_readdata_pre_23;
input 	av_readdata_pre_11;
input 	av_readdata_pre_13;
input 	av_readdata_pre_161;
input 	av_readdata_pre_12;
input 	av_readdata_pre_14;
input 	av_readdata_pre_15;
input 	av_readdata_pre_181;
input 	av_readdata_pre_171;
input 	av_readdata_pre_10;
input 	av_readdata_pre_9;
input 	av_readdata_pre_8;
input 	av_readdata_pre_211;
input 	av_readdata_pre_191;
input 	av_readdata_pre_201;
input 	av_readdata_pre_81;
input 	av_readdata_pre_82;
output 	src_data_8;
input 	av_readdata_pre_121;
input 	av_readdata_pre_122;
output 	src_data_12;
input 	av_readdata_pre_111;
output 	src_data_11;
input 	av_readdata_pre_101;
input 	av_readdata_pre_102;
output 	src_data_10;
input 	av_readdata_pre_91;
input 	av_readdata_pre_92;
output 	src_data_9;
input 	av_readdata_pre_151;
input 	av_readdata_pre_152;
output 	src_data_15;
input 	av_readdata_pre_141;
input 	av_readdata_pre_142;
output 	src_data_14;
input 	av_readdata_pre_131;
input 	av_readdata_pre_132;
output 	src_data_13;
input 	av_readdata_pre_162;
output 	src_data_16;
input 	av_readdata_pre_202;
output 	src_data_20;
input 	av_readdata_pre_192;
output 	src_data_19;
input 	av_readdata_pre_182;
output 	src_data_18;
input 	av_readdata_pre_172;
output 	src_data_17;
input 	av_readdata_pre_231;
output 	src_data_23;
input 	av_readdata_pre_222;
output 	src_data_22;
input 	av_readdata_pre_212;
output 	src_data_21;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \src_payload~0_combout ;
wire \src_data[8]~0_combout ;
wire \src_payload~1_combout ;
wire \src_data[12]~2_combout ;
wire \src_data[11]~4_combout ;
wire \src_payload~2_combout ;
wire \src_data[10]~5_combout ;
wire \src_payload~3_combout ;
wire \src_data[9]~7_combout ;
wire \src_payload~4_combout ;
wire \src_data[15]~9_combout ;
wire \src_payload~5_combout ;
wire \src_data[14]~11_combout ;
wire \src_payload~6_combout ;
wire \src_data[13]~13_combout ;
wire \src_payload~7_combout ;
wire \src_data[16]~15_combout ;
wire \src_payload~8_combout ;
wire \src_data[20]~17_combout ;
wire \src_payload~9_combout ;
wire \src_data[19]~19_combout ;
wire \src_payload~10_combout ;
wire \src_data[18]~21_combout ;
wire \src_payload~11_combout ;
wire \src_data[17]~23_combout ;
wire \src_data[23]~25_combout ;
wire \src_payload~12_combout ;
wire \src_data[22]~26_combout ;
wire \src_payload~13_combout ;
wire \src_data[21]~28_combout ;


cycloneive_lcell_comb \WideOr1~0 (
	.dataa(mem_73_0),
	.datab(mem_55_0),
	.datac(read_latency_shift_reg_01),
	.datad(read_latency_shift_reg_02),
	.cin(gnd),
	.combout(WideOr11),
	.cout());
defparam \WideOr1~0 .lut_mask = 16'hEFFF;
defparam \WideOr1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb WideOr1(
	.dataa(WideOr11),
	.datab(read_latency_shift_reg_0),
	.datac(read_latency_shift_reg_03),
	.datad(read_latency_shift_reg_04),
	.cin(gnd),
	.combout(WideOr12),
	.cout());
defparam WideOr1.lut_mask = 16'hBFFF;
defparam WideOr1.sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr1~1 (
	.dataa(gnd),
	.datab(read_latency_shift_reg_0),
	.datac(read_latency_shift_reg_03),
	.datad(read_latency_shift_reg_04),
	.cin(gnd),
	.combout(WideOr13),
	.cout());
defparam \WideOr1~1 .lut_mask = 16'h3FFF;
defparam \WideOr1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[8]~1 (
	.dataa(\src_payload~0_combout ),
	.datab(\src_data[8]~0_combout ),
	.datac(read_latency_shift_reg_04),
	.datad(q_b_8),
	.cin(gnd),
	.combout(src_data_8),
	.cout());
defparam \src_data[8]~1 .lut_mask = 16'hFFFE;
defparam \src_data[8]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[12]~3 (
	.dataa(\src_payload~1_combout ),
	.datab(\src_data[12]~2_combout ),
	.datac(read_latency_shift_reg_04),
	.datad(q_b_12),
	.cin(gnd),
	.combout(src_data_12),
	.cout());
defparam \src_data[12]~3 .lut_mask = 16'hFFFE;
defparam \src_data[12]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[11] (
	.dataa(\src_data[11]~4_combout ),
	.datab(src0_valid),
	.datac(av_readdata_pre_11),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_11),
	.cout());
defparam \src_data[11] .lut_mask = 16'hFEFE;
defparam \src_data[11] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[10]~6 (
	.dataa(\src_payload~2_combout ),
	.datab(\src_data[10]~5_combout ),
	.datac(read_latency_shift_reg_04),
	.datad(q_b_10),
	.cin(gnd),
	.combout(src_data_10),
	.cout());
defparam \src_data[10]~6 .lut_mask = 16'hFFFE;
defparam \src_data[10]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[9]~8 (
	.dataa(\src_payload~3_combout ),
	.datab(\src_data[9]~7_combout ),
	.datac(read_latency_shift_reg_04),
	.datad(q_b_9),
	.cin(gnd),
	.combout(src_data_9),
	.cout());
defparam \src_data[9]~8 .lut_mask = 16'hFFFE;
defparam \src_data[9]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[15]~10 (
	.dataa(\src_payload~4_combout ),
	.datab(\src_data[15]~9_combout ),
	.datac(read_latency_shift_reg_04),
	.datad(q_b_15),
	.cin(gnd),
	.combout(src_data_15),
	.cout());
defparam \src_data[15]~10 .lut_mask = 16'hFFFE;
defparam \src_data[15]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[14]~12 (
	.dataa(\src_payload~5_combout ),
	.datab(\src_data[14]~11_combout ),
	.datac(read_latency_shift_reg_04),
	.datad(q_b_14),
	.cin(gnd),
	.combout(src_data_14),
	.cout());
defparam \src_data[14]~12 .lut_mask = 16'hFFFE;
defparam \src_data[14]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[13]~14 (
	.dataa(\src_payload~6_combout ),
	.datab(\src_data[13]~13_combout ),
	.datac(read_latency_shift_reg_04),
	.datad(q_b_13),
	.cin(gnd),
	.combout(src_data_13),
	.cout());
defparam \src_data[13]~14 .lut_mask = 16'hFFFE;
defparam \src_data[13]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[16]~16 (
	.dataa(\src_payload~7_combout ),
	.datab(\src_data[16]~15_combout ),
	.datac(read_latency_shift_reg_04),
	.datad(q_b_16),
	.cin(gnd),
	.combout(src_data_16),
	.cout());
defparam \src_data[16]~16 .lut_mask = 16'hFFFE;
defparam \src_data[16]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[20]~18 (
	.dataa(\src_payload~8_combout ),
	.datab(\src_data[20]~17_combout ),
	.datac(read_latency_shift_reg_04),
	.datad(q_b_20),
	.cin(gnd),
	.combout(src_data_20),
	.cout());
defparam \src_data[20]~18 .lut_mask = 16'hFFFE;
defparam \src_data[20]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[19]~20 (
	.dataa(\src_payload~9_combout ),
	.datab(\src_data[19]~19_combout ),
	.datac(read_latency_shift_reg_04),
	.datad(q_b_19),
	.cin(gnd),
	.combout(src_data_19),
	.cout());
defparam \src_data[19]~20 .lut_mask = 16'hFFFE;
defparam \src_data[19]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[18]~22 (
	.dataa(\src_payload~10_combout ),
	.datab(\src_data[18]~21_combout ),
	.datac(read_latency_shift_reg_04),
	.datad(q_b_18),
	.cin(gnd),
	.combout(src_data_18),
	.cout());
defparam \src_data[18]~22 .lut_mask = 16'hFFFE;
defparam \src_data[18]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[17]~24 (
	.dataa(\src_payload~11_combout ),
	.datab(\src_data[17]~23_combout ),
	.datac(read_latency_shift_reg_04),
	.datad(q_b_17),
	.cin(gnd),
	.combout(src_data_17),
	.cout());
defparam \src_data[17]~24 .lut_mask = 16'hFFFE;
defparam \src_data[17]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[23] (
	.dataa(\src_data[23]~25_combout ),
	.datab(src0_valid),
	.datac(av_readdata_pre_23),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_23),
	.cout());
defparam \src_data[23] .lut_mask = 16'hFEFE;
defparam \src_data[23] .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[22]~27 (
	.dataa(\src_payload~12_combout ),
	.datab(\src_data[22]~26_combout ),
	.datac(read_latency_shift_reg_04),
	.datad(q_b_22),
	.cin(gnd),
	.combout(src_data_22),
	.cout());
defparam \src_data[22]~27 .lut_mask = 16'hFFFE;
defparam \src_data[22]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[21]~29 (
	.dataa(\src_payload~13_combout ),
	.datab(\src_data[21]~28_combout ),
	.datac(read_latency_shift_reg_04),
	.datad(q_b_21),
	.cin(gnd),
	.combout(src_data_21),
	.cout());
defparam \src_data[21]~29 .lut_mask = 16'hFFFE;
defparam \src_data[21]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~0 (
	.dataa(read_latency_shift_reg_01),
	.datab(av_readdata_pre_8),
	.datac(mem_73_0),
	.datad(mem_55_0),
	.cin(gnd),
	.combout(\src_payload~0_combout ),
	.cout());
defparam \src_payload~0 .lut_mask = 16'hEFFF;
defparam \src_payload~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[8]~0 (
	.dataa(read_latency_shift_reg_02),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_81),
	.datad(av_readdata_pre_82),
	.cin(gnd),
	.combout(\src_data[8]~0_combout ),
	.cout());
defparam \src_data[8]~0 .lut_mask = 16'hFFFE;
defparam \src_data[8]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~1 (
	.dataa(read_latency_shift_reg_01),
	.datab(av_readdata_pre_12),
	.datac(mem_73_0),
	.datad(mem_55_0),
	.cin(gnd),
	.combout(\src_payload~1_combout ),
	.cout());
defparam \src_payload~1 .lut_mask = 16'hEFFF;
defparam \src_payload~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[12]~2 (
	.dataa(read_latency_shift_reg_02),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_121),
	.datad(av_readdata_pre_122),
	.cin(gnd),
	.combout(\src_data[12]~2_combout ),
	.cout());
defparam \src_data[12]~2 .lut_mask = 16'hFFFE;
defparam \src_data[12]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[11]~4 (
	.dataa(read_latency_shift_reg_03),
	.datab(read_latency_shift_reg_04),
	.datac(q_b_11),
	.datad(av_readdata_pre_111),
	.cin(gnd),
	.combout(\src_data[11]~4_combout ),
	.cout());
defparam \src_data[11]~4 .lut_mask = 16'hFFFE;
defparam \src_data[11]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~2 (
	.dataa(read_latency_shift_reg_01),
	.datab(av_readdata_pre_10),
	.datac(mem_73_0),
	.datad(mem_55_0),
	.cin(gnd),
	.combout(\src_payload~2_combout ),
	.cout());
defparam \src_payload~2 .lut_mask = 16'hEFFF;
defparam \src_payload~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[10]~5 (
	.dataa(read_latency_shift_reg_02),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_101),
	.datad(av_readdata_pre_102),
	.cin(gnd),
	.combout(\src_data[10]~5_combout ),
	.cout());
defparam \src_data[10]~5 .lut_mask = 16'hFFFE;
defparam \src_data[10]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~3 (
	.dataa(read_latency_shift_reg_01),
	.datab(av_readdata_pre_9),
	.datac(mem_73_0),
	.datad(mem_55_0),
	.cin(gnd),
	.combout(\src_payload~3_combout ),
	.cout());
defparam \src_payload~3 .lut_mask = 16'hEFFF;
defparam \src_payload~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[9]~7 (
	.dataa(read_latency_shift_reg_02),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_91),
	.datad(av_readdata_pre_92),
	.cin(gnd),
	.combout(\src_data[9]~7_combout ),
	.cout());
defparam \src_data[9]~7 .lut_mask = 16'hFFFE;
defparam \src_data[9]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~4 (
	.dataa(read_latency_shift_reg_01),
	.datab(av_readdata_pre_15),
	.datac(mem_73_0),
	.datad(mem_55_0),
	.cin(gnd),
	.combout(\src_payload~4_combout ),
	.cout());
defparam \src_payload~4 .lut_mask = 16'hEFFF;
defparam \src_payload~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[15]~9 (
	.dataa(read_latency_shift_reg_02),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_151),
	.datad(av_readdata_pre_152),
	.cin(gnd),
	.combout(\src_data[15]~9_combout ),
	.cout());
defparam \src_data[15]~9 .lut_mask = 16'hFFFE;
defparam \src_data[15]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~5 (
	.dataa(read_latency_shift_reg_01),
	.datab(av_readdata_pre_14),
	.datac(mem_73_0),
	.datad(mem_55_0),
	.cin(gnd),
	.combout(\src_payload~5_combout ),
	.cout());
defparam \src_payload~5 .lut_mask = 16'hEFFF;
defparam \src_payload~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[14]~11 (
	.dataa(read_latency_shift_reg_02),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_141),
	.datad(av_readdata_pre_142),
	.cin(gnd),
	.combout(\src_data[14]~11_combout ),
	.cout());
defparam \src_data[14]~11 .lut_mask = 16'hFFFE;
defparam \src_data[14]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~6 (
	.dataa(read_latency_shift_reg_01),
	.datab(av_readdata_pre_13),
	.datac(mem_73_0),
	.datad(mem_55_0),
	.cin(gnd),
	.combout(\src_payload~6_combout ),
	.cout());
defparam \src_payload~6 .lut_mask = 16'hEFFF;
defparam \src_payload~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[13]~13 (
	.dataa(read_latency_shift_reg_02),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_131),
	.datad(av_readdata_pre_132),
	.cin(gnd),
	.combout(\src_data[13]~13_combout ),
	.cout());
defparam \src_data[13]~13 .lut_mask = 16'hFFFE;
defparam \src_data[13]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~7 (
	.dataa(read_latency_shift_reg_01),
	.datab(av_readdata_pre_161),
	.datac(mem_73_0),
	.datad(mem_55_0),
	.cin(gnd),
	.combout(\src_payload~7_combout ),
	.cout());
defparam \src_payload~7 .lut_mask = 16'hEFFF;
defparam \src_payload~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[16]~15 (
	.dataa(read_latency_shift_reg_02),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_162),
	.datad(av_readdata_pre_16),
	.cin(gnd),
	.combout(\src_data[16]~15_combout ),
	.cout());
defparam \src_data[16]~15 .lut_mask = 16'hFFFE;
defparam \src_data[16]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~8 (
	.dataa(read_latency_shift_reg_01),
	.datab(av_readdata_pre_201),
	.datac(mem_73_0),
	.datad(mem_55_0),
	.cin(gnd),
	.combout(\src_payload~8_combout ),
	.cout());
defparam \src_payload~8 .lut_mask = 16'hEFFF;
defparam \src_payload~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[20]~17 (
	.dataa(read_latency_shift_reg_02),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_202),
	.datad(av_readdata_pre_20),
	.cin(gnd),
	.combout(\src_data[20]~17_combout ),
	.cout());
defparam \src_data[20]~17 .lut_mask = 16'hFFFE;
defparam \src_data[20]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~9 (
	.dataa(read_latency_shift_reg_01),
	.datab(av_readdata_pre_191),
	.datac(mem_73_0),
	.datad(mem_55_0),
	.cin(gnd),
	.combout(\src_payload~9_combout ),
	.cout());
defparam \src_payload~9 .lut_mask = 16'hEFFF;
defparam \src_payload~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[19]~19 (
	.dataa(read_latency_shift_reg_02),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_192),
	.datad(av_readdata_pre_19),
	.cin(gnd),
	.combout(\src_data[19]~19_combout ),
	.cout());
defparam \src_data[19]~19 .lut_mask = 16'hFFFE;
defparam \src_data[19]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~10 (
	.dataa(read_latency_shift_reg_01),
	.datab(av_readdata_pre_181),
	.datac(mem_73_0),
	.datad(mem_55_0),
	.cin(gnd),
	.combout(\src_payload~10_combout ),
	.cout());
defparam \src_payload~10 .lut_mask = 16'hEFFF;
defparam \src_payload~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[18]~21 (
	.dataa(read_latency_shift_reg_02),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_182),
	.datad(av_readdata_pre_18),
	.cin(gnd),
	.combout(\src_data[18]~21_combout ),
	.cout());
defparam \src_data[18]~21 .lut_mask = 16'hFFFE;
defparam \src_data[18]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~11 (
	.dataa(read_latency_shift_reg_01),
	.datab(av_readdata_pre_171),
	.datac(mem_73_0),
	.datad(mem_55_0),
	.cin(gnd),
	.combout(\src_payload~11_combout ),
	.cout());
defparam \src_payload~11 .lut_mask = 16'hEFFF;
defparam \src_payload~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[17]~23 (
	.dataa(read_latency_shift_reg_02),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_172),
	.datad(av_readdata_pre_17),
	.cin(gnd),
	.combout(\src_data[17]~23_combout ),
	.cout());
defparam \src_data[17]~23 .lut_mask = 16'hFFFE;
defparam \src_data[17]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[23]~25 (
	.dataa(read_latency_shift_reg_03),
	.datab(read_latency_shift_reg_04),
	.datac(q_b_23),
	.datad(av_readdata_pre_231),
	.cin(gnd),
	.combout(\src_data[23]~25_combout ),
	.cout());
defparam \src_data[23]~25 .lut_mask = 16'hFFFE;
defparam \src_data[23]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~12 (
	.dataa(read_latency_shift_reg_01),
	.datab(av_readdata_pre_221),
	.datac(mem_73_0),
	.datad(mem_55_0),
	.cin(gnd),
	.combout(\src_payload~12_combout ),
	.cout());
defparam \src_payload~12 .lut_mask = 16'hEFFF;
defparam \src_payload~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[22]~26 (
	.dataa(read_latency_shift_reg_02),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_222),
	.datad(av_readdata_pre_22),
	.cin(gnd),
	.combout(\src_data[22]~26_combout ),
	.cout());
defparam \src_data[22]~26 .lut_mask = 16'hFFFE;
defparam \src_data[22]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~13 (
	.dataa(read_latency_shift_reg_01),
	.datab(av_readdata_pre_211),
	.datac(mem_73_0),
	.datad(mem_55_0),
	.cin(gnd),
	.combout(\src_payload~13_combout ),
	.cout());
defparam \src_payload~13 .lut_mask = 16'hEFFF;
defparam \src_payload~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[21]~28 (
	.dataa(read_latency_shift_reg_02),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_212),
	.datad(av_readdata_pre_21),
	.cin(gnd),
	.combout(\src_data[21]~28_combout ),
	.cout());
defparam \src_data[21]~28 .lut_mask = 16'hFFFE;
defparam \src_data[21]~28 .sum_lutc_input = "datac";

endmodule

module nios_mcu_nios_mcu_mm_interconnect_0_rsp_mux_001 (
	q_a_11,
	q_a_13,
	q_a_16,
	q_a_1,
	q_a_3,
	q_a_5,
	q_a_4,
	q_a_15,
	q_a_21,
	q_a_19,
	q_a_20,
	read_latency_shift_reg_0,
	src_payload,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10)/* synthesis synthesis_greybox=1 */;
input 	q_a_11;
input 	q_a_13;
input 	q_a_16;
input 	q_a_1;
input 	q_a_3;
input 	q_a_5;
input 	q_a_4;
input 	q_a_15;
input 	q_a_21;
input 	q_a_19;
input 	q_a_20;
input 	read_latency_shift_reg_0;
output 	src_payload;
output 	src_payload1;
output 	src_payload2;
output 	src_payload3;
output 	src_payload4;
output 	src_payload5;
output 	src_payload6;
output 	src_payload7;
output 	src_payload8;
output 	src_payload9;
output 	src_payload10;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \src_payload~0 (
	.dataa(read_latency_shift_reg_0),
	.datab(q_a_11),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload),
	.cout());
defparam \src_payload~0 .lut_mask = 16'hEEEE;
defparam \src_payload~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~1 (
	.dataa(read_latency_shift_reg_0),
	.datab(q_a_13),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload1),
	.cout());
defparam \src_payload~1 .lut_mask = 16'hEEEE;
defparam \src_payload~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~2 (
	.dataa(read_latency_shift_reg_0),
	.datab(q_a_16),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload2),
	.cout());
defparam \src_payload~2 .lut_mask = 16'hEEEE;
defparam \src_payload~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~3 (
	.dataa(read_latency_shift_reg_0),
	.datab(q_a_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload3),
	.cout());
defparam \src_payload~3 .lut_mask = 16'hEEEE;
defparam \src_payload~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~4 (
	.dataa(read_latency_shift_reg_0),
	.datab(q_a_3),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload4),
	.cout());
defparam \src_payload~4 .lut_mask = 16'hEEEE;
defparam \src_payload~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~5 (
	.dataa(read_latency_shift_reg_0),
	.datab(q_a_5),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload5),
	.cout());
defparam \src_payload~5 .lut_mask = 16'hEEEE;
defparam \src_payload~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~6 (
	.dataa(read_latency_shift_reg_0),
	.datab(q_a_4),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload6),
	.cout());
defparam \src_payload~6 .lut_mask = 16'hEEEE;
defparam \src_payload~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~7 (
	.dataa(read_latency_shift_reg_0),
	.datab(q_a_15),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload7),
	.cout());
defparam \src_payload~7 .lut_mask = 16'hEEEE;
defparam \src_payload~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~8 (
	.dataa(read_latency_shift_reg_0),
	.datab(q_a_21),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload8),
	.cout());
defparam \src_payload~8 .lut_mask = 16'hEEEE;
defparam \src_payload~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~9 (
	.dataa(read_latency_shift_reg_0),
	.datab(q_a_19),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload9),
	.cout());
defparam \src_payload~9 .lut_mask = 16'hEEEE;
defparam \src_payload~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~10 (
	.dataa(read_latency_shift_reg_0),
	.datab(q_a_20),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload10),
	.cout());
defparam \src_payload~10 .lut_mask = 16'hEEEE;
defparam \src_payload~10 .sum_lutc_input = "datac";

endmodule

module nios_mcu_nios_mcu_nios_cpu (
	sr_0,
	W_alu_result_12,
	W_alu_result_15,
	W_alu_result_14,
	W_alu_result_13,
	W_alu_result_11,
	W_alu_result_10,
	W_alu_result_9,
	W_alu_result_8,
	W_alu_result_7,
	W_alu_result_6,
	W_alu_result_5,
	W_alu_result_4,
	W_alu_result_3,
	W_alu_result_2,
	q_a_0,
	q_b_0,
	q_a_22,
	q_a_23,
	q_a_24,
	q_b_24,
	q_a_25,
	q_b_25,
	q_a_26,
	q_b_26,
	q_a_12,
	q_b_1,
	q_b_3,
	q_a_2,
	q_b_2,
	q_b_5,
	q_b_4,
	q_a_14,
	q_a_18,
	q_a_17,
	q_a_10,
	q_a_9,
	q_a_8,
	q_a_7,
	q_b_7,
	q_a_6,
	q_b_6,
	readdata_0,
	d_writedata_24,
	d_writedata_25,
	d_writedata_26,
	readdata_1,
	readdata_3,
	readdata_2,
	q_a_27,
	q_b_27,
	q_a_28,
	q_b_28,
	q_a_29,
	q_b_29,
	q_a_30,
	q_b_30,
	q_a_31,
	q_b_31,
	d_writedata_27,
	d_writedata_28,
	d_writedata_29,
	d_writedata_30,
	d_writedata_31,
	ir_out_0,
	ir_out_1,
	d_writedata_0,
	r_sync_rst,
	d_write,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	read_latency_shift_reg_0,
	d_read,
	m0_write,
	mem_73_0,
	mem_55_0,
	read_latency_shift_reg_01,
	read_latency_shift_reg_02,
	WideOr1,
	read_latency_shift_reg_03,
	read_latency_shift_reg_04,
	WideOr11,
	saved_grant_0,
	debug_mem_slave_waitrequest,
	mem_used_1,
	av_waitrequest,
	F_pc_10,
	F_pc_9,
	F_pc_8,
	F_pc_7,
	F_pc_6,
	F_pc_5,
	F_pc_4,
	F_pc_3,
	F_pc_2,
	F_pc_1,
	F_pc_0,
	F_pc_13,
	F_pc_12,
	F_pc_11,
	i_read,
	WideOr12,
	rf_source_valid,
	hbreak_enabled,
	WideOr13,
	av_readdata_pre_0,
	av_readdata_pre_01,
	av_readdata_pre_02,
	src0_valid,
	av_readdata_pre_03,
	av_readdata_pre_22,
	read_latency_shift_reg_05,
	src1_valid,
	av_readdata_pre_23,
	av_readdata_pre_24,
	av_readdata_pre_25,
	av_readdata_pre_26,
	src_payload,
	av_readdata_pre_11,
	src_payload1,
	av_readdata_pre_13,
	src_payload2,
	av_readdata_pre_16,
	av_readdata_pre_12,
	src_payload3,
	av_readdata_pre_1,
	src_payload4,
	av_readdata_pre_3,
	av_readdata_pre_2,
	src_payload5,
	av_readdata_pre_5,
	src_payload6,
	av_readdata_pre_4,
	av_readdata_pre_14,
	src_payload7,
	av_readdata_pre_15,
	av_readdata_pre_18,
	av_readdata_pre_17,
	av_readdata_pre_10,
	av_readdata_pre_9,
	av_readdata_pre_8,
	av_readdata_pre_7,
	av_readdata_pre_6,
	src_payload8,
	av_readdata_pre_21,
	src_payload9,
	av_readdata_pre_19,
	src_payload10,
	av_readdata_pre_20,
	src_data_46,
	av_readdata_pre_110,
	av_readdata_pre_111,
	av_readdata_pre_112,
	av_readdata_pre_27,
	av_readdata_pre_28,
	av_readdata_pre_29,
	av_readdata_pre_31,
	av_readdata_pre_32,
	av_readdata_pre_33,
	av_readdata_pre_41,
	av_readdata_pre_42,
	av_readdata_pre_43,
	av_readdata_pre_51,
	av_readdata_pre_52,
	av_readdata_pre_53,
	av_readdata_pre_61,
	av_readdata_pre_62,
	av_readdata_pre_63,
	av_readdata_pre_71,
	av_readdata_pre_72,
	av_readdata_pre_73,
	r_early_rst,
	src_data_8,
	d_byteenable_0,
	av_readdata_9,
	av_readdata_8,
	readdata_22,
	d_writedata_22,
	d_byteenable_2,
	readdata_23,
	d_writedata_23,
	readdata_24,
	d_byteenable_3,
	readdata_25,
	readdata_26,
	d_writedata_11,
	d_byteenable_1,
	readdata_11,
	d_writedata_13,
	readdata_13,
	d_writedata_16,
	readdata_16,
	readdata_12,
	d_writedata_12,
	readdata_5,
	readdata_4,
	d_writedata_14,
	readdata_14,
	d_writedata_15,
	readdata_15,
	d_writedata_18,
	readdata_18,
	src_data_12,
	av_readdata_pre_271,
	av_readdata_pre_281,
	av_readdata_pre_291,
	av_readdata_pre_30,
	av_readdata_pre_311,
	d_writedata_17,
	readdata_17,
	src_data_11,
	src_data_10,
	src_data_9,
	readdata_10,
	d_writedata_10,
	readdata_9,
	d_writedata_9,
	readdata_8,
	d_writedata_8,
	readdata_7,
	readdata_6,
	d_writedata_21,
	readdata_21,
	src_data_15,
	d_writedata_19,
	readdata_19,
	d_writedata_20,
	readdata_20,
	src_data_14,
	src_data_13,
	src_payload11,
	src_payload12,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_32,
	src_data_16,
	src_data_20,
	readdata_27,
	readdata_28,
	readdata_29,
	readdata_30,
	readdata_31,
	src_data_19,
	src_data_18,
	src_data_17,
	src_data_23,
	src_data_22,
	src_data_21,
	src_payload13,
	av_readdata_pre_241,
	av_readdata_pre_312,
	av_readdata_pre_301,
	av_readdata_pre_292,
	av_readdata_pre_282,
	av_readdata_pre_272,
	av_readdata_pre_261,
	av_readdata_pre_251,
	src_payload14,
	src_payload15,
	src_payload16,
	src_data_34,
	src_payload17,
	src_payload18,
	src_data_35,
	src_payload19,
	src_payload20,
	src_payload21,
	src_data_33,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32,
	src_payload33,
	src_payload34,
	src_payload35,
	src_payload36,
	src_payload37,
	src_payload38,
	src_payload39,
	src_payload40,
	src_payload41,
	src_payload42,
	src_payload43,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	sr_0;
output 	W_alu_result_12;
output 	W_alu_result_15;
output 	W_alu_result_14;
output 	W_alu_result_13;
output 	W_alu_result_11;
output 	W_alu_result_10;
output 	W_alu_result_9;
output 	W_alu_result_8;
output 	W_alu_result_7;
output 	W_alu_result_6;
output 	W_alu_result_5;
output 	W_alu_result_4;
output 	W_alu_result_3;
output 	W_alu_result_2;
input 	q_a_0;
input 	q_b_0;
input 	q_a_22;
input 	q_a_23;
input 	q_a_24;
input 	q_b_24;
input 	q_a_25;
input 	q_b_25;
input 	q_a_26;
input 	q_b_26;
input 	q_a_12;
input 	q_b_1;
input 	q_b_3;
input 	q_a_2;
input 	q_b_2;
input 	q_b_5;
input 	q_b_4;
input 	q_a_14;
input 	q_a_18;
input 	q_a_17;
input 	q_a_10;
input 	q_a_9;
input 	q_a_8;
input 	q_a_7;
input 	q_b_7;
input 	q_a_6;
input 	q_b_6;
output 	readdata_0;
output 	d_writedata_24;
output 	d_writedata_25;
output 	d_writedata_26;
output 	readdata_1;
output 	readdata_3;
output 	readdata_2;
input 	q_a_27;
input 	q_b_27;
input 	q_a_28;
input 	q_b_28;
input 	q_a_29;
input 	q_b_29;
input 	q_a_30;
input 	q_b_30;
input 	q_a_31;
input 	q_b_31;
output 	d_writedata_27;
output 	d_writedata_28;
output 	d_writedata_29;
output 	d_writedata_30;
output 	d_writedata_31;
output 	ir_out_0;
output 	ir_out_1;
output 	d_writedata_0;
input 	r_sync_rst;
output 	d_write;
output 	d_writedata_1;
output 	d_writedata_2;
output 	d_writedata_3;
output 	d_writedata_4;
output 	d_writedata_5;
output 	d_writedata_6;
output 	d_writedata_7;
input 	read_latency_shift_reg_0;
output 	d_read;
input 	m0_write;
input 	mem_73_0;
input 	mem_55_0;
input 	read_latency_shift_reg_01;
input 	read_latency_shift_reg_02;
input 	WideOr1;
input 	read_latency_shift_reg_03;
input 	read_latency_shift_reg_04;
input 	WideOr11;
input 	saved_grant_0;
output 	debug_mem_slave_waitrequest;
input 	mem_used_1;
input 	av_waitrequest;
output 	F_pc_10;
output 	F_pc_9;
output 	F_pc_8;
output 	F_pc_7;
output 	F_pc_6;
output 	F_pc_5;
output 	F_pc_4;
output 	F_pc_3;
output 	F_pc_2;
output 	F_pc_1;
output 	F_pc_0;
output 	F_pc_13;
output 	F_pc_12;
output 	F_pc_11;
output 	i_read;
input 	WideOr12;
input 	rf_source_valid;
output 	hbreak_enabled;
input 	WideOr13;
input 	av_readdata_pre_0;
input 	av_readdata_pre_01;
input 	av_readdata_pre_02;
input 	src0_valid;
input 	av_readdata_pre_03;
input 	av_readdata_pre_22;
input 	read_latency_shift_reg_05;
input 	src1_valid;
input 	av_readdata_pre_23;
input 	av_readdata_pre_24;
input 	av_readdata_pre_25;
input 	av_readdata_pre_26;
input 	src_payload;
input 	av_readdata_pre_11;
input 	src_payload1;
input 	av_readdata_pre_13;
input 	src_payload2;
input 	av_readdata_pre_16;
input 	av_readdata_pre_12;
input 	src_payload3;
input 	av_readdata_pre_1;
input 	src_payload4;
input 	av_readdata_pre_3;
input 	av_readdata_pre_2;
input 	src_payload5;
input 	av_readdata_pre_5;
input 	src_payload6;
input 	av_readdata_pre_4;
input 	av_readdata_pre_14;
input 	src_payload7;
input 	av_readdata_pre_15;
input 	av_readdata_pre_18;
input 	av_readdata_pre_17;
input 	av_readdata_pre_10;
input 	av_readdata_pre_9;
input 	av_readdata_pre_8;
input 	av_readdata_pre_7;
input 	av_readdata_pre_6;
input 	src_payload8;
input 	av_readdata_pre_21;
input 	src_payload9;
input 	av_readdata_pre_19;
input 	src_payload10;
input 	av_readdata_pre_20;
input 	src_data_46;
input 	av_readdata_pre_110;
input 	av_readdata_pre_111;
input 	av_readdata_pre_112;
input 	av_readdata_pre_27;
input 	av_readdata_pre_28;
input 	av_readdata_pre_29;
input 	av_readdata_pre_31;
input 	av_readdata_pre_32;
input 	av_readdata_pre_33;
input 	av_readdata_pre_41;
input 	av_readdata_pre_42;
input 	av_readdata_pre_43;
input 	av_readdata_pre_51;
input 	av_readdata_pre_52;
input 	av_readdata_pre_53;
input 	av_readdata_pre_61;
input 	av_readdata_pre_62;
input 	av_readdata_pre_63;
input 	av_readdata_pre_71;
input 	av_readdata_pre_72;
input 	av_readdata_pre_73;
input 	r_early_rst;
input 	src_data_8;
output 	d_byteenable_0;
input 	av_readdata_9;
input 	av_readdata_8;
output 	readdata_22;
output 	d_writedata_22;
output 	d_byteenable_2;
output 	readdata_23;
output 	d_writedata_23;
output 	readdata_24;
output 	d_byteenable_3;
output 	readdata_25;
output 	readdata_26;
output 	d_writedata_11;
output 	d_byteenable_1;
output 	readdata_11;
output 	d_writedata_13;
output 	readdata_13;
output 	d_writedata_16;
output 	readdata_16;
output 	readdata_12;
output 	d_writedata_12;
output 	readdata_5;
output 	readdata_4;
output 	d_writedata_14;
output 	readdata_14;
output 	d_writedata_15;
output 	readdata_15;
output 	d_writedata_18;
output 	readdata_18;
input 	src_data_12;
input 	av_readdata_pre_271;
input 	av_readdata_pre_281;
input 	av_readdata_pre_291;
input 	av_readdata_pre_30;
input 	av_readdata_pre_311;
output 	d_writedata_17;
output 	readdata_17;
input 	src_data_11;
input 	src_data_10;
input 	src_data_9;
output 	readdata_10;
output 	d_writedata_10;
output 	readdata_9;
output 	d_writedata_9;
output 	readdata_8;
output 	d_writedata_8;
output 	readdata_7;
output 	readdata_6;
output 	d_writedata_21;
output 	readdata_21;
input 	src_data_15;
output 	d_writedata_19;
output 	readdata_19;
output 	d_writedata_20;
output 	readdata_20;
input 	src_data_14;
input 	src_data_13;
input 	src_payload11;
input 	src_payload12;
input 	src_data_38;
input 	src_data_39;
input 	src_data_40;
input 	src_data_41;
input 	src_data_42;
input 	src_data_43;
input 	src_data_44;
input 	src_data_45;
input 	src_data_32;
input 	src_data_16;
input 	src_data_20;
output 	readdata_27;
output 	readdata_28;
output 	readdata_29;
output 	readdata_30;
output 	readdata_31;
input 	src_data_19;
input 	src_data_18;
input 	src_data_17;
input 	src_data_23;
input 	src_data_22;
input 	src_data_21;
input 	src_payload13;
input 	av_readdata_pre_241;
input 	av_readdata_pre_312;
input 	av_readdata_pre_301;
input 	av_readdata_pre_292;
input 	av_readdata_pre_282;
input 	av_readdata_pre_272;
input 	av_readdata_pre_261;
input 	av_readdata_pre_251;
input 	src_payload14;
input 	src_payload15;
input 	src_payload16;
input 	src_data_34;
input 	src_payload17;
input 	src_payload18;
input 	src_data_35;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_data_33;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	src_payload32;
input 	src_payload33;
input 	src_payload34;
input 	src_payload35;
input 	src_payload36;
input 	src_payload37;
input 	src_payload38;
input 	src_payload39;
input 	src_payload40;
input 	src_payload41;
input 	src_payload42;
input 	src_payload43;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nios_mcu_nios_mcu_nios_cpu_cpu cpu(
	.sr_0(sr_0),
	.W_alu_result_12(W_alu_result_12),
	.W_alu_result_15(W_alu_result_15),
	.W_alu_result_14(W_alu_result_14),
	.W_alu_result_13(W_alu_result_13),
	.W_alu_result_11(W_alu_result_11),
	.W_alu_result_10(W_alu_result_10),
	.W_alu_result_9(W_alu_result_9),
	.W_alu_result_8(W_alu_result_8),
	.W_alu_result_7(W_alu_result_7),
	.W_alu_result_6(W_alu_result_6),
	.W_alu_result_5(W_alu_result_5),
	.W_alu_result_4(W_alu_result_4),
	.W_alu_result_3(W_alu_result_3),
	.W_alu_result_2(W_alu_result_2),
	.q_a_0(q_a_0),
	.q_b_0(q_b_0),
	.q_a_22(q_a_22),
	.q_a_23(q_a_23),
	.q_a_24(q_a_24),
	.q_b_24(q_b_24),
	.q_a_25(q_a_25),
	.q_b_25(q_b_25),
	.q_a_26(q_a_26),
	.q_b_26(q_b_26),
	.q_a_12(q_a_12),
	.q_b_1(q_b_1),
	.q_b_3(q_b_3),
	.q_a_2(q_a_2),
	.q_b_2(q_b_2),
	.q_b_5(q_b_5),
	.q_b_4(q_b_4),
	.q_a_14(q_a_14),
	.q_a_18(q_a_18),
	.q_a_17(q_a_17),
	.q_a_10(q_a_10),
	.q_a_9(q_a_9),
	.q_a_8(q_a_8),
	.q_a_7(q_a_7),
	.q_b_7(q_b_7),
	.q_a_6(q_a_6),
	.q_b_6(q_b_6),
	.readdata_0(readdata_0),
	.d_writedata_24(d_writedata_24),
	.d_writedata_25(d_writedata_25),
	.d_writedata_26(d_writedata_26),
	.readdata_1(readdata_1),
	.readdata_3(readdata_3),
	.readdata_2(readdata_2),
	.q_a_27(q_a_27),
	.q_b_27(q_b_27),
	.q_a_28(q_a_28),
	.q_b_28(q_b_28),
	.q_a_29(q_a_29),
	.q_b_29(q_b_29),
	.q_a_30(q_a_30),
	.q_b_30(q_b_30),
	.q_a_31(q_a_31),
	.q_b_31(q_b_31),
	.d_writedata_27(d_writedata_27),
	.d_writedata_28(d_writedata_28),
	.d_writedata_29(d_writedata_29),
	.d_writedata_30(d_writedata_30),
	.d_writedata_31(d_writedata_31),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.d_writedata_0(d_writedata_0),
	.r_sync_rst(r_sync_rst),
	.d_write1(d_write),
	.d_writedata_1(d_writedata_1),
	.d_writedata_2(d_writedata_2),
	.d_writedata_3(d_writedata_3),
	.d_writedata_4(d_writedata_4),
	.d_writedata_5(d_writedata_5),
	.d_writedata_6(d_writedata_6),
	.d_writedata_7(d_writedata_7),
	.read_latency_shift_reg_0(read_latency_shift_reg_0),
	.d_read1(d_read),
	.m0_write(m0_write),
	.mem_73_0(mem_73_0),
	.mem_55_0(mem_55_0),
	.read_latency_shift_reg_01(read_latency_shift_reg_01),
	.read_latency_shift_reg_02(read_latency_shift_reg_02),
	.WideOr1(WideOr1),
	.read_latency_shift_reg_03(read_latency_shift_reg_03),
	.read_latency_shift_reg_04(read_latency_shift_reg_04),
	.WideOr11(WideOr11),
	.saved_grant_0(saved_grant_0),
	.debug_mem_slave_waitrequest(debug_mem_slave_waitrequest),
	.mem_used_1(mem_used_1),
	.av_waitrequest(av_waitrequest),
	.F_pc_10(F_pc_10),
	.F_pc_9(F_pc_9),
	.F_pc_8(F_pc_8),
	.F_pc_7(F_pc_7),
	.F_pc_6(F_pc_6),
	.F_pc_5(F_pc_5),
	.F_pc_4(F_pc_4),
	.F_pc_3(F_pc_3),
	.F_pc_2(F_pc_2),
	.F_pc_1(F_pc_1),
	.F_pc_0(F_pc_0),
	.F_pc_13(F_pc_13),
	.F_pc_12(F_pc_12),
	.F_pc_11(F_pc_11),
	.i_read1(i_read),
	.WideOr12(WideOr12),
	.rf_source_valid(rf_source_valid),
	.hbreak_enabled1(hbreak_enabled),
	.WideOr13(WideOr13),
	.av_readdata_pre_0(av_readdata_pre_0),
	.av_readdata_pre_01(av_readdata_pre_01),
	.av_readdata_pre_02(av_readdata_pre_02),
	.src0_valid(src0_valid),
	.av_readdata_pre_03(av_readdata_pre_03),
	.av_readdata_pre_22(av_readdata_pre_22),
	.read_latency_shift_reg_05(read_latency_shift_reg_05),
	.src1_valid(src1_valid),
	.av_readdata_pre_23(av_readdata_pre_23),
	.av_readdata_pre_24(av_readdata_pre_24),
	.av_readdata_pre_25(av_readdata_pre_25),
	.av_readdata_pre_26(av_readdata_pre_26),
	.src_payload(src_payload),
	.av_readdata_pre_11(av_readdata_pre_11),
	.src_payload1(src_payload1),
	.av_readdata_pre_13(av_readdata_pre_13),
	.src_payload2(src_payload2),
	.av_readdata_pre_16(av_readdata_pre_16),
	.av_readdata_pre_12(av_readdata_pre_12),
	.src_payload3(src_payload3),
	.av_readdata_pre_1(av_readdata_pre_1),
	.src_payload4(src_payload4),
	.av_readdata_pre_3(av_readdata_pre_3),
	.av_readdata_pre_2(av_readdata_pre_2),
	.src_payload5(src_payload5),
	.av_readdata_pre_5(av_readdata_pre_5),
	.src_payload6(src_payload6),
	.av_readdata_pre_4(av_readdata_pre_4),
	.av_readdata_pre_14(av_readdata_pre_14),
	.src_payload7(src_payload7),
	.av_readdata_pre_15(av_readdata_pre_15),
	.av_readdata_pre_18(av_readdata_pre_18),
	.av_readdata_pre_17(av_readdata_pre_17),
	.av_readdata_pre_10(av_readdata_pre_10),
	.av_readdata_pre_9(av_readdata_pre_9),
	.av_readdata_pre_8(av_readdata_pre_8),
	.av_readdata_pre_7(av_readdata_pre_7),
	.av_readdata_pre_6(av_readdata_pre_6),
	.src_payload8(src_payload8),
	.av_readdata_pre_21(av_readdata_pre_21),
	.src_payload9(src_payload9),
	.av_readdata_pre_19(av_readdata_pre_19),
	.src_payload10(src_payload10),
	.av_readdata_pre_20(av_readdata_pre_20),
	.src_data_46(src_data_46),
	.av_readdata_pre_110(av_readdata_pre_110),
	.av_readdata_pre_111(av_readdata_pre_111),
	.av_readdata_pre_112(av_readdata_pre_112),
	.av_readdata_pre_27(av_readdata_pre_27),
	.av_readdata_pre_28(av_readdata_pre_28),
	.av_readdata_pre_29(av_readdata_pre_29),
	.av_readdata_pre_31(av_readdata_pre_31),
	.av_readdata_pre_32(av_readdata_pre_32),
	.av_readdata_pre_33(av_readdata_pre_33),
	.av_readdata_pre_41(av_readdata_pre_41),
	.av_readdata_pre_42(av_readdata_pre_42),
	.av_readdata_pre_43(av_readdata_pre_43),
	.av_readdata_pre_51(av_readdata_pre_51),
	.av_readdata_pre_52(av_readdata_pre_52),
	.av_readdata_pre_53(av_readdata_pre_53),
	.av_readdata_pre_61(av_readdata_pre_61),
	.av_readdata_pre_62(av_readdata_pre_62),
	.av_readdata_pre_63(av_readdata_pre_63),
	.av_readdata_pre_71(av_readdata_pre_71),
	.av_readdata_pre_72(av_readdata_pre_72),
	.av_readdata_pre_73(av_readdata_pre_73),
	.r_early_rst(r_early_rst),
	.src_data_8(src_data_8),
	.d_byteenable_0(d_byteenable_0),
	.av_readdata_9(av_readdata_9),
	.av_readdata_8(av_readdata_8),
	.readdata_22(readdata_22),
	.d_writedata_22(d_writedata_22),
	.d_byteenable_2(d_byteenable_2),
	.readdata_23(readdata_23),
	.d_writedata_23(d_writedata_23),
	.readdata_24(readdata_24),
	.d_byteenable_3(d_byteenable_3),
	.readdata_25(readdata_25),
	.readdata_26(readdata_26),
	.d_writedata_11(d_writedata_11),
	.d_byteenable_1(d_byteenable_1),
	.readdata_11(readdata_11),
	.d_writedata_13(d_writedata_13),
	.readdata_13(readdata_13),
	.d_writedata_16(d_writedata_16),
	.readdata_16(readdata_16),
	.readdata_12(readdata_12),
	.d_writedata_12(d_writedata_12),
	.readdata_5(readdata_5),
	.readdata_4(readdata_4),
	.d_writedata_14(d_writedata_14),
	.readdata_14(readdata_14),
	.d_writedata_15(d_writedata_15),
	.readdata_15(readdata_15),
	.d_writedata_18(d_writedata_18),
	.readdata_18(readdata_18),
	.src_data_12(src_data_12),
	.av_readdata_pre_271(av_readdata_pre_271),
	.av_readdata_pre_281(av_readdata_pre_281),
	.av_readdata_pre_291(av_readdata_pre_291),
	.av_readdata_pre_30(av_readdata_pre_30),
	.av_readdata_pre_311(av_readdata_pre_311),
	.d_writedata_17(d_writedata_17),
	.readdata_17(readdata_17),
	.src_data_11(src_data_11),
	.src_data_10(src_data_10),
	.src_data_9(src_data_9),
	.readdata_10(readdata_10),
	.d_writedata_10(d_writedata_10),
	.readdata_9(readdata_9),
	.d_writedata_9(d_writedata_9),
	.readdata_8(readdata_8),
	.d_writedata_8(d_writedata_8),
	.readdata_7(readdata_7),
	.readdata_6(readdata_6),
	.d_writedata_21(d_writedata_21),
	.readdata_21(readdata_21),
	.src_data_15(src_data_15),
	.d_writedata_19(d_writedata_19),
	.readdata_19(readdata_19),
	.d_writedata_20(d_writedata_20),
	.readdata_20(readdata_20),
	.src_data_14(src_data_14),
	.src_data_13(src_data_13),
	.src_payload11(src_payload11),
	.src_payload12(src_payload12),
	.src_data_38(src_data_38),
	.src_data_39(src_data_39),
	.src_data_40(src_data_40),
	.src_data_41(src_data_41),
	.src_data_42(src_data_42),
	.src_data_43(src_data_43),
	.src_data_44(src_data_44),
	.src_data_45(src_data_45),
	.src_data_32(src_data_32),
	.src_data_16(src_data_16),
	.src_data_20(src_data_20),
	.readdata_27(readdata_27),
	.readdata_28(readdata_28),
	.readdata_29(readdata_29),
	.readdata_30(readdata_30),
	.readdata_31(readdata_31),
	.src_data_19(src_data_19),
	.src_data_18(src_data_18),
	.src_data_17(src_data_17),
	.src_data_23(src_data_23),
	.src_data_22(src_data_22),
	.src_data_21(src_data_21),
	.src_payload13(src_payload13),
	.av_readdata_pre_241(av_readdata_pre_241),
	.av_readdata_pre_312(av_readdata_pre_312),
	.av_readdata_pre_301(av_readdata_pre_301),
	.av_readdata_pre_292(av_readdata_pre_292),
	.av_readdata_pre_282(av_readdata_pre_282),
	.av_readdata_pre_272(av_readdata_pre_272),
	.av_readdata_pre_261(av_readdata_pre_261),
	.av_readdata_pre_251(av_readdata_pre_251),
	.src_payload14(src_payload14),
	.src_payload15(src_payload15),
	.src_payload16(src_payload16),
	.src_data_34(src_data_34),
	.src_payload17(src_payload17),
	.src_payload18(src_payload18),
	.src_data_35(src_data_35),
	.src_payload19(src_payload19),
	.src_payload20(src_payload20),
	.src_payload21(src_payload21),
	.src_data_33(src_data_33),
	.src_payload22(src_payload22),
	.src_payload23(src_payload23),
	.src_payload24(src_payload24),
	.src_payload25(src_payload25),
	.src_payload26(src_payload26),
	.src_payload27(src_payload27),
	.src_payload28(src_payload28),
	.src_payload29(src_payload29),
	.src_payload30(src_payload30),
	.src_payload31(src_payload31),
	.src_payload32(src_payload32),
	.src_payload33(src_payload33),
	.src_payload34(src_payload34),
	.src_payload35(src_payload35),
	.src_payload36(src_payload36),
	.src_payload37(src_payload37),
	.src_payload38(src_payload38),
	.src_payload39(src_payload39),
	.src_payload40(src_payload40),
	.src_payload41(src_payload41),
	.src_payload42(src_payload42),
	.src_payload43(src_payload43),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_1(state_1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3),
	.irf_reg_0_2(irf_reg_0_2),
	.irf_reg_1_2(irf_reg_1_2),
	.clk_clk(clk_clk));

endmodule

module nios_mcu_nios_mcu_nios_cpu_cpu (
	sr_0,
	W_alu_result_12,
	W_alu_result_15,
	W_alu_result_14,
	W_alu_result_13,
	W_alu_result_11,
	W_alu_result_10,
	W_alu_result_9,
	W_alu_result_8,
	W_alu_result_7,
	W_alu_result_6,
	W_alu_result_5,
	W_alu_result_4,
	W_alu_result_3,
	W_alu_result_2,
	q_a_0,
	q_b_0,
	q_a_22,
	q_a_23,
	q_a_24,
	q_b_24,
	q_a_25,
	q_b_25,
	q_a_26,
	q_b_26,
	q_a_12,
	q_b_1,
	q_b_3,
	q_a_2,
	q_b_2,
	q_b_5,
	q_b_4,
	q_a_14,
	q_a_18,
	q_a_17,
	q_a_10,
	q_a_9,
	q_a_8,
	q_a_7,
	q_b_7,
	q_a_6,
	q_b_6,
	readdata_0,
	d_writedata_24,
	d_writedata_25,
	d_writedata_26,
	readdata_1,
	readdata_3,
	readdata_2,
	q_a_27,
	q_b_27,
	q_a_28,
	q_b_28,
	q_a_29,
	q_b_29,
	q_a_30,
	q_b_30,
	q_a_31,
	q_b_31,
	d_writedata_27,
	d_writedata_28,
	d_writedata_29,
	d_writedata_30,
	d_writedata_31,
	ir_out_0,
	ir_out_1,
	d_writedata_0,
	r_sync_rst,
	d_write1,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	read_latency_shift_reg_0,
	d_read1,
	m0_write,
	mem_73_0,
	mem_55_0,
	read_latency_shift_reg_01,
	read_latency_shift_reg_02,
	WideOr1,
	read_latency_shift_reg_03,
	read_latency_shift_reg_04,
	WideOr11,
	saved_grant_0,
	debug_mem_slave_waitrequest,
	mem_used_1,
	av_waitrequest,
	F_pc_10,
	F_pc_9,
	F_pc_8,
	F_pc_7,
	F_pc_6,
	F_pc_5,
	F_pc_4,
	F_pc_3,
	F_pc_2,
	F_pc_1,
	F_pc_0,
	F_pc_13,
	F_pc_12,
	F_pc_11,
	i_read1,
	WideOr12,
	rf_source_valid,
	hbreak_enabled1,
	WideOr13,
	av_readdata_pre_0,
	av_readdata_pre_01,
	av_readdata_pre_02,
	src0_valid,
	av_readdata_pre_03,
	av_readdata_pre_22,
	read_latency_shift_reg_05,
	src1_valid,
	av_readdata_pre_23,
	av_readdata_pre_24,
	av_readdata_pre_25,
	av_readdata_pre_26,
	src_payload,
	av_readdata_pre_11,
	src_payload1,
	av_readdata_pre_13,
	src_payload2,
	av_readdata_pre_16,
	av_readdata_pre_12,
	src_payload3,
	av_readdata_pre_1,
	src_payload4,
	av_readdata_pre_3,
	av_readdata_pre_2,
	src_payload5,
	av_readdata_pre_5,
	src_payload6,
	av_readdata_pre_4,
	av_readdata_pre_14,
	src_payload7,
	av_readdata_pre_15,
	av_readdata_pre_18,
	av_readdata_pre_17,
	av_readdata_pre_10,
	av_readdata_pre_9,
	av_readdata_pre_8,
	av_readdata_pre_7,
	av_readdata_pre_6,
	src_payload8,
	av_readdata_pre_21,
	src_payload9,
	av_readdata_pre_19,
	src_payload10,
	av_readdata_pre_20,
	src_data_46,
	av_readdata_pre_110,
	av_readdata_pre_111,
	av_readdata_pre_112,
	av_readdata_pre_27,
	av_readdata_pre_28,
	av_readdata_pre_29,
	av_readdata_pre_31,
	av_readdata_pre_32,
	av_readdata_pre_33,
	av_readdata_pre_41,
	av_readdata_pre_42,
	av_readdata_pre_43,
	av_readdata_pre_51,
	av_readdata_pre_52,
	av_readdata_pre_53,
	av_readdata_pre_61,
	av_readdata_pre_62,
	av_readdata_pre_63,
	av_readdata_pre_71,
	av_readdata_pre_72,
	av_readdata_pre_73,
	r_early_rst,
	src_data_8,
	d_byteenable_0,
	av_readdata_9,
	av_readdata_8,
	readdata_22,
	d_writedata_22,
	d_byteenable_2,
	readdata_23,
	d_writedata_23,
	readdata_24,
	d_byteenable_3,
	readdata_25,
	readdata_26,
	d_writedata_11,
	d_byteenable_1,
	readdata_11,
	d_writedata_13,
	readdata_13,
	d_writedata_16,
	readdata_16,
	readdata_12,
	d_writedata_12,
	readdata_5,
	readdata_4,
	d_writedata_14,
	readdata_14,
	d_writedata_15,
	readdata_15,
	d_writedata_18,
	readdata_18,
	src_data_12,
	av_readdata_pre_271,
	av_readdata_pre_281,
	av_readdata_pre_291,
	av_readdata_pre_30,
	av_readdata_pre_311,
	d_writedata_17,
	readdata_17,
	src_data_11,
	src_data_10,
	src_data_9,
	readdata_10,
	d_writedata_10,
	readdata_9,
	d_writedata_9,
	readdata_8,
	d_writedata_8,
	readdata_7,
	readdata_6,
	d_writedata_21,
	readdata_21,
	src_data_15,
	d_writedata_19,
	readdata_19,
	d_writedata_20,
	readdata_20,
	src_data_14,
	src_data_13,
	src_payload11,
	src_payload12,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_32,
	src_data_16,
	src_data_20,
	readdata_27,
	readdata_28,
	readdata_29,
	readdata_30,
	readdata_31,
	src_data_19,
	src_data_18,
	src_data_17,
	src_data_23,
	src_data_22,
	src_data_21,
	src_payload13,
	av_readdata_pre_241,
	av_readdata_pre_312,
	av_readdata_pre_301,
	av_readdata_pre_292,
	av_readdata_pre_282,
	av_readdata_pre_272,
	av_readdata_pre_261,
	av_readdata_pre_251,
	src_payload14,
	src_payload15,
	src_payload16,
	src_data_34,
	src_payload17,
	src_payload18,
	src_data_35,
	src_payload19,
	src_payload20,
	src_payload21,
	src_data_33,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32,
	src_payload33,
	src_payload34,
	src_payload35,
	src_payload36,
	src_payload37,
	src_payload38,
	src_payload39,
	src_payload40,
	src_payload41,
	src_payload42,
	src_payload43,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	sr_0;
output 	W_alu_result_12;
output 	W_alu_result_15;
output 	W_alu_result_14;
output 	W_alu_result_13;
output 	W_alu_result_11;
output 	W_alu_result_10;
output 	W_alu_result_9;
output 	W_alu_result_8;
output 	W_alu_result_7;
output 	W_alu_result_6;
output 	W_alu_result_5;
output 	W_alu_result_4;
output 	W_alu_result_3;
output 	W_alu_result_2;
input 	q_a_0;
input 	q_b_0;
input 	q_a_22;
input 	q_a_23;
input 	q_a_24;
input 	q_b_24;
input 	q_a_25;
input 	q_b_25;
input 	q_a_26;
input 	q_b_26;
input 	q_a_12;
input 	q_b_1;
input 	q_b_3;
input 	q_a_2;
input 	q_b_2;
input 	q_b_5;
input 	q_b_4;
input 	q_a_14;
input 	q_a_18;
input 	q_a_17;
input 	q_a_10;
input 	q_a_9;
input 	q_a_8;
input 	q_a_7;
input 	q_b_7;
input 	q_a_6;
input 	q_b_6;
output 	readdata_0;
output 	d_writedata_24;
output 	d_writedata_25;
output 	d_writedata_26;
output 	readdata_1;
output 	readdata_3;
output 	readdata_2;
input 	q_a_27;
input 	q_b_27;
input 	q_a_28;
input 	q_b_28;
input 	q_a_29;
input 	q_b_29;
input 	q_a_30;
input 	q_b_30;
input 	q_a_31;
input 	q_b_31;
output 	d_writedata_27;
output 	d_writedata_28;
output 	d_writedata_29;
output 	d_writedata_30;
output 	d_writedata_31;
output 	ir_out_0;
output 	ir_out_1;
output 	d_writedata_0;
input 	r_sync_rst;
output 	d_write1;
output 	d_writedata_1;
output 	d_writedata_2;
output 	d_writedata_3;
output 	d_writedata_4;
output 	d_writedata_5;
output 	d_writedata_6;
output 	d_writedata_7;
input 	read_latency_shift_reg_0;
output 	d_read1;
input 	m0_write;
input 	mem_73_0;
input 	mem_55_0;
input 	read_latency_shift_reg_01;
input 	read_latency_shift_reg_02;
input 	WideOr1;
input 	read_latency_shift_reg_03;
input 	read_latency_shift_reg_04;
input 	WideOr11;
input 	saved_grant_0;
output 	debug_mem_slave_waitrequest;
input 	mem_used_1;
input 	av_waitrequest;
output 	F_pc_10;
output 	F_pc_9;
output 	F_pc_8;
output 	F_pc_7;
output 	F_pc_6;
output 	F_pc_5;
output 	F_pc_4;
output 	F_pc_3;
output 	F_pc_2;
output 	F_pc_1;
output 	F_pc_0;
output 	F_pc_13;
output 	F_pc_12;
output 	F_pc_11;
output 	i_read1;
input 	WideOr12;
input 	rf_source_valid;
output 	hbreak_enabled1;
input 	WideOr13;
input 	av_readdata_pre_0;
input 	av_readdata_pre_01;
input 	av_readdata_pre_02;
input 	src0_valid;
input 	av_readdata_pre_03;
input 	av_readdata_pre_22;
input 	read_latency_shift_reg_05;
input 	src1_valid;
input 	av_readdata_pre_23;
input 	av_readdata_pre_24;
input 	av_readdata_pre_25;
input 	av_readdata_pre_26;
input 	src_payload;
input 	av_readdata_pre_11;
input 	src_payload1;
input 	av_readdata_pre_13;
input 	src_payload2;
input 	av_readdata_pre_16;
input 	av_readdata_pre_12;
input 	src_payload3;
input 	av_readdata_pre_1;
input 	src_payload4;
input 	av_readdata_pre_3;
input 	av_readdata_pre_2;
input 	src_payload5;
input 	av_readdata_pre_5;
input 	src_payload6;
input 	av_readdata_pre_4;
input 	av_readdata_pre_14;
input 	src_payload7;
input 	av_readdata_pre_15;
input 	av_readdata_pre_18;
input 	av_readdata_pre_17;
input 	av_readdata_pre_10;
input 	av_readdata_pre_9;
input 	av_readdata_pre_8;
input 	av_readdata_pre_7;
input 	av_readdata_pre_6;
input 	src_payload8;
input 	av_readdata_pre_21;
input 	src_payload9;
input 	av_readdata_pre_19;
input 	src_payload10;
input 	av_readdata_pre_20;
input 	src_data_46;
input 	av_readdata_pre_110;
input 	av_readdata_pre_111;
input 	av_readdata_pre_112;
input 	av_readdata_pre_27;
input 	av_readdata_pre_28;
input 	av_readdata_pre_29;
input 	av_readdata_pre_31;
input 	av_readdata_pre_32;
input 	av_readdata_pre_33;
input 	av_readdata_pre_41;
input 	av_readdata_pre_42;
input 	av_readdata_pre_43;
input 	av_readdata_pre_51;
input 	av_readdata_pre_52;
input 	av_readdata_pre_53;
input 	av_readdata_pre_61;
input 	av_readdata_pre_62;
input 	av_readdata_pre_63;
input 	av_readdata_pre_71;
input 	av_readdata_pre_72;
input 	av_readdata_pre_73;
input 	r_early_rst;
input 	src_data_8;
output 	d_byteenable_0;
input 	av_readdata_9;
input 	av_readdata_8;
output 	readdata_22;
output 	d_writedata_22;
output 	d_byteenable_2;
output 	readdata_23;
output 	d_writedata_23;
output 	readdata_24;
output 	d_byteenable_3;
output 	readdata_25;
output 	readdata_26;
output 	d_writedata_11;
output 	d_byteenable_1;
output 	readdata_11;
output 	d_writedata_13;
output 	readdata_13;
output 	d_writedata_16;
output 	readdata_16;
output 	readdata_12;
output 	d_writedata_12;
output 	readdata_5;
output 	readdata_4;
output 	d_writedata_14;
output 	readdata_14;
output 	d_writedata_15;
output 	readdata_15;
output 	d_writedata_18;
output 	readdata_18;
input 	src_data_12;
input 	av_readdata_pre_271;
input 	av_readdata_pre_281;
input 	av_readdata_pre_291;
input 	av_readdata_pre_30;
input 	av_readdata_pre_311;
output 	d_writedata_17;
output 	readdata_17;
input 	src_data_11;
input 	src_data_10;
input 	src_data_9;
output 	readdata_10;
output 	d_writedata_10;
output 	readdata_9;
output 	d_writedata_9;
output 	readdata_8;
output 	d_writedata_8;
output 	readdata_7;
output 	readdata_6;
output 	d_writedata_21;
output 	readdata_21;
input 	src_data_15;
output 	d_writedata_19;
output 	readdata_19;
output 	d_writedata_20;
output 	readdata_20;
input 	src_data_14;
input 	src_data_13;
input 	src_payload11;
input 	src_payload12;
input 	src_data_38;
input 	src_data_39;
input 	src_data_40;
input 	src_data_41;
input 	src_data_42;
input 	src_data_43;
input 	src_data_44;
input 	src_data_45;
input 	src_data_32;
input 	src_data_16;
input 	src_data_20;
output 	readdata_27;
output 	readdata_28;
output 	readdata_29;
output 	readdata_30;
output 	readdata_31;
input 	src_data_19;
input 	src_data_18;
input 	src_data_17;
input 	src_data_23;
input 	src_data_22;
input 	src_data_21;
input 	src_payload13;
input 	av_readdata_pre_241;
input 	av_readdata_pre_312;
input 	av_readdata_pre_301;
input 	av_readdata_pre_292;
input 	av_readdata_pre_282;
input 	av_readdata_pre_272;
input 	av_readdata_pre_261;
input 	av_readdata_pre_251;
input 	src_payload14;
input 	src_payload15;
input 	src_payload16;
input 	src_data_34;
input 	src_payload17;
input 	src_payload18;
input 	src_data_35;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_data_33;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	src_payload32;
input 	src_payload33;
input 	src_payload34;
input 	src_payload35;
input 	src_payload36;
input 	src_payload37;
input 	src_payload38;
input 	src_payload39;
input 	src_payload40;
input 	src_payload41;
input 	src_payload42;
input 	src_payload43;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ;
wire \W_alu_result[0]~q ;
wire \nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[12] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[11] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[10] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[9] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[8] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[7] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[6] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[5] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[4] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[3] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[2] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[1] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[0] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[15] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[14] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[13] ;
wire \W_alu_result[1]~q ;
wire \av_ld_byte1_data[0]~q ;
wire \Add1~66_combout ;
wire \Add1~68_combout ;
wire \Add1~70_combout ;
wire \Add1~72_combout ;
wire \Add1~74_combout ;
wire \Add1~76_combout ;
wire \Add1~78_combout ;
wire \Add1~80_combout ;
wire \Add1~82_combout ;
wire \Add1~84_combout ;
wire \Add1~86_combout ;
wire \Add1~88_combout ;
wire \Add1~90_combout ;
wire \Add1~92_combout ;
wire \Add1~94_combout ;
wire \Add1~96_combout ;
wire \W_alu_result[0]~14_combout ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci|the_nios_mcu_nios_cpu_cpu_nios2_oci_debug|jtag_break~q ;
wire \av_ld_byte1_data[4]~q ;
wire \av_ld_byte1_data[3]~q ;
wire \av_ld_byte1_data[2]~q ;
wire \av_ld_byte1_data[1]~q ;
wire \av_ld_byte1_data[7]~q ;
wire \av_ld_byte1_data[6]~q ;
wire \av_ld_byte1_data[5]~q ;
wire \W_alu_result[1]~15_combout ;
wire \av_ld_byte1_data[0]~0_combout ;
wire \av_ld_byte2_data[0]~q ;
wire \nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[31] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[31] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[16] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[16] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[30] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[30] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[29] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[29] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[28] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[28] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[27] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[27] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[26] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[26] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[25] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[25] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[24] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[24] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[23] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[23] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[22] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[22] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[21] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[21] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[20] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[20] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[19] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[19] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[18] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[18] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[17] ;
wire \nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[17] ;
wire \av_ld_byte1_data[4]~4_combout ;
wire \av_ld_byte2_data[4]~q ;
wire \av_ld_byte1_data[3]~5_combout ;
wire \av_ld_byte2_data[3]~q ;
wire \av_ld_byte1_data[2]~6_combout ;
wire \av_ld_byte2_data[2]~q ;
wire \av_ld_byte1_data[1]~7_combout ;
wire \av_ld_byte2_data[1]~q ;
wire \av_ld_byte1_data[7]~1_combout ;
wire \av_ld_byte2_data[7]~q ;
wire \av_ld_byte1_data[6]~2_combout ;
wire \av_ld_byte2_data[6]~q ;
wire \av_ld_byte1_data[5]~3_combout ;
wire \av_ld_byte2_data[5]~q ;
wire \av_ld_byte2_data[0]~0_combout ;
wire \W_alu_result[31]~q ;
wire \W_alu_result[16]~q ;
wire \W_alu_result[30]~q ;
wire \W_alu_result[29]~q ;
wire \W_alu_result[28]~q ;
wire \W_alu_result[27]~q ;
wire \W_alu_result[26]~q ;
wire \W_alu_result[25]~q ;
wire \W_alu_result[24]~q ;
wire \W_alu_result[23]~q ;
wire \W_alu_result[22]~q ;
wire \W_alu_result[21]~q ;
wire \W_alu_result[20]~q ;
wire \W_alu_result[19]~q ;
wire \W_alu_result[18]~q ;
wire \W_alu_result[17]~q ;
wire \av_ld_byte2_data[4]~4_combout ;
wire \av_ld_byte2_data[3]~5_combout ;
wire \av_ld_byte2_data[2]~6_combout ;
wire \av_ld_byte2_data[1]~7_combout ;
wire \av_ld_byte2_data[7]~1_combout ;
wire \av_ld_byte2_data[6]~2_combout ;
wire \av_ld_byte2_data[5]~3_combout ;
wire \W_alu_result[31]~16_combout ;
wire \W_alu_result[16]~17_combout ;
wire \W_alu_result[30]~18_combout ;
wire \W_alu_result[29]~19_combout ;
wire \W_alu_result[28]~20_combout ;
wire \W_alu_result[27]~21_combout ;
wire \W_alu_result[26]~22_combout ;
wire \W_alu_result[25]~23_combout ;
wire \W_alu_result[24]~24_combout ;
wire \W_alu_result[23]~25_combout ;
wire \W_alu_result[22]~26_combout ;
wire \W_alu_result[21]~27_combout ;
wire \W_alu_result[20]~28_combout ;
wire \W_alu_result[19]~29_combout ;
wire \W_alu_result[18]~30_combout ;
wire \W_alu_result[17]~31_combout ;
wire \R_wr_dst_reg~q ;
wire \W_rf_wren~combout ;
wire \av_ld_byte0_data[0]~q ;
wire \W_rf_wr_data[0]~0_combout ;
wire \W_control_rd_data[0]~q ;
wire \W_rf_wr_data[0]~1_combout ;
wire \W_rf_wr_data[0]~2_combout ;
wire \R_dst_regnum[0]~q ;
wire \R_dst_regnum[1]~q ;
wire \R_dst_regnum[2]~q ;
wire \R_dst_regnum[3]~q ;
wire \R_dst_regnum[4]~q ;
wire \D_iw[22]~q ;
wire \D_iw[23]~q ;
wire \D_iw[24]~q ;
wire \D_iw[25]~q ;
wire \D_iw[26]~q ;
wire \av_ld_byte0_data[1]~q ;
wire \W_rf_wr_data[1]~3_combout ;
wire \av_ld_byte0_data[2]~q ;
wire \W_rf_wr_data[2]~4_combout ;
wire \av_ld_byte0_data[3]~q ;
wire \W_rf_wr_data[3]~5_combout ;
wire \av_ld_byte0_data[4]~q ;
wire \W_rf_wr_data[4]~6_combout ;
wire \av_ld_byte0_data[5]~q ;
wire \W_rf_wr_data[5]~7_combout ;
wire \av_ld_byte0_data[6]~q ;
wire \W_rf_wr_data[6]~8_combout ;
wire \av_ld_byte0_data[7]~q ;
wire \W_rf_wr_data[7]~9_combout ;
wire \D_wr_dst_reg~0_combout ;
wire \D_wr_dst_reg~1_combout ;
wire \Equal0~14_combout ;
wire \D_ctrl_implicit_dst_eretaddr~14_combout ;
wire \D_ctrl_implicit_dst_eretaddr~15_combout ;
wire \D_ctrl_implicit_dst_eretaddr~17_combout ;
wire \D_dst_regnum[1]~0_combout ;
wire \D_dst_regnum[1]~1_combout ;
wire \D_dst_regnum[4]~2_combout ;
wire \D_dst_regnum[4]~3_combout ;
wire \D_dst_regnum[3]~4_combout ;
wire \D_dst_regnum[3]~5_combout ;
wire \D_dst_regnum[4]~6_combout ;
wire \D_dst_regnum[4]~7_combout ;
wire \D_dst_regnum[2]~8_combout ;
wire \Equal0~18_combout ;
wire \D_dst_regnum[0]~9_combout ;
wire \D_wr_dst_reg~2_combout ;
wire \av_ld_byte0_data_nxt[0]~16_combout ;
wire \av_ld_byte0_data_nxt[0]~17_combout ;
wire \av_ld_byte0_data_nxt[0]~18_combout ;
wire \av_ld_rshift8~0_combout ;
wire \av_ld_rshift8~1_combout ;
wire \av_ld_byte0_data[7]~0_combout ;
wire \E_control_rd_data[0]~0_combout ;
wire \E_control_rd_data[0]~1_combout ;
wire \E_control_rd_data[0]~2_combout ;
wire \E_control_rd_data[0]~3_combout ;
wire \D_ctrl_ld_signed~1_combout ;
wire \F_iw[22]~0_combout ;
wire \F_iw[22]~1_combout ;
wire \F_iw[23]~2_combout ;
wire \F_iw[23]~3_combout ;
wire \F_iw[24]~4_combout ;
wire \F_iw[24]~5_combout ;
wire \F_iw[25]~6_combout ;
wire \F_iw[25]~7_combout ;
wire \F_iw[26]~8_combout ;
wire \F_iw[26]~9_combout ;
wire \W_rf_wr_data[12]~10_combout ;
wire \D_iw[27]~q ;
wire \D_iw[28]~q ;
wire \D_iw[29]~q ;
wire \D_iw[30]~q ;
wire \D_iw[31]~q ;
wire \W_rf_wr_data[11]~11_combout ;
wire \W_rf_wr_data[10]~12_combout ;
wire \W_rf_wr_data[9]~13_combout ;
wire \W_rf_wr_data[8]~14_combout ;
wire \W_rf_wr_data[15]~15_combout ;
wire \W_rf_wr_data[14]~16_combout ;
wire \W_rf_wr_data[13]~17_combout ;
wire \av_ld_byte0_data_nxt[1]~19_combout ;
wire \av_ld_byte0_data_nxt[1]~20_combout ;
wire \av_ld_byte0_data_nxt[1]~21_combout ;
wire \av_ld_byte0_data_nxt[2]~22_combout ;
wire \av_ld_byte0_data_nxt[2]~23_combout ;
wire \av_ld_byte0_data_nxt[2]~24_combout ;
wire \av_ld_byte0_data_nxt[3]~25_combout ;
wire \av_ld_byte0_data_nxt[3]~26_combout ;
wire \av_ld_byte0_data_nxt[3]~27_combout ;
wire \av_ld_byte0_data_nxt[4]~28_combout ;
wire \av_ld_byte0_data_nxt[4]~29_combout ;
wire \av_ld_byte0_data_nxt[4]~30_combout ;
wire \av_ld_byte0_data_nxt[5]~31_combout ;
wire \av_ld_byte0_data_nxt[5]~32_combout ;
wire \av_ld_byte0_data_nxt[5]~33_combout ;
wire \av_ld_byte0_data_nxt[6]~34_combout ;
wire \av_ld_byte0_data_nxt[6]~35_combout ;
wire \av_ld_byte0_data_nxt[6]~36_combout ;
wire \av_ld_byte0_data_nxt[7]~37_combout ;
wire \av_ld_byte0_data_nxt[7]~38_combout ;
wire \av_ld_byte0_data_nxt[7]~39_combout ;
wire \R_ctrl_ld_signed~q ;
wire \av_fill_bit~0_combout ;
wire \av_ld_byte1_data_en~0_combout ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci|the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_ienable[0]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci|the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_single_step_mode~q ;
wire \F_iw[27]~43_combout ;
wire \F_iw[27]~44_combout ;
wire \F_iw[28]~45_combout ;
wire \F_iw[28]~46_combout ;
wire \F_iw[29]~47_combout ;
wire \F_iw[29]~48_combout ;
wire \F_iw[30]~49_combout ;
wire \F_iw[30]~50_combout ;
wire \F_iw[31]~51_combout ;
wire \F_iw[31]~52_combout ;
wire \av_ld_byte3_data[0]~q ;
wire \av_ld_byte3_data[7]~q ;
wire \W_rf_wr_data[31]~18_combout ;
wire \W_rf_wr_data[16]~19_combout ;
wire \av_ld_byte3_data[6]~q ;
wire \W_rf_wr_data[30]~20_combout ;
wire \av_ld_byte3_data[5]~q ;
wire \W_rf_wr_data[29]~21_combout ;
wire \av_ld_byte3_data[4]~q ;
wire \W_rf_wr_data[28]~22_combout ;
wire \av_ld_byte3_data[3]~q ;
wire \W_rf_wr_data[27]~23_combout ;
wire \av_ld_byte3_data[2]~q ;
wire \W_rf_wr_data[26]~24_combout ;
wire \av_ld_byte3_data[1]~q ;
wire \W_rf_wr_data[25]~25_combout ;
wire \W_rf_wr_data[24]~26_combout ;
wire \W_rf_wr_data[23]~27_combout ;
wire \W_rf_wr_data[22]~28_combout ;
wire \W_rf_wr_data[21]~29_combout ;
wire \W_rf_wr_data[20]~30_combout ;
wire \W_rf_wr_data[19]~31_combout ;
wire \W_rf_wr_data[18]~32_combout ;
wire \W_rf_wr_data[17]~33_combout ;
wire \av_ld_byte3_data_nxt~0_combout ;
wire \av_ld_byte3_data_nxt~1_combout ;
wire \av_ld_byte3_data_nxt~2_combout ;
wire \av_ld_byte3_data_nxt~3_combout ;
wire \av_ld_byte3_data_nxt~4_combout ;
wire \av_ld_byte3_data_nxt~5_combout ;
wire \av_ld_byte3_data_nxt~6_combout ;
wire \av_ld_byte3_data_nxt~7_combout ;
wire \av_ld_byte3_data_nxt~8_combout ;
wire \av_ld_byte3_data_nxt~9_combout ;
wire \av_ld_byte3_data_nxt~10_combout ;
wire \av_ld_byte3_data_nxt~11_combout ;
wire \av_ld_byte3_data_nxt~12_combout ;
wire \av_ld_byte3_data_nxt~13_combout ;
wire \av_ld_byte3_data_nxt~14_combout ;
wire \av_ld_byte3_data_nxt~15_combout ;
wire \av_ld_byte3_data_nxt~16_combout ;
wire \av_ld_byte3_data_nxt~17_combout ;
wire \av_ld_byte3_data_nxt~18_combout ;
wire \av_ld_byte3_data_nxt~19_combout ;
wire \av_ld_byte3_data_nxt~20_combout ;
wire \av_ld_byte3_data_nxt~21_combout ;
wire \av_ld_byte3_data_nxt~22_combout ;
wire \av_ld_byte3_data_nxt~23_combout ;
wire \av_ld_byte0_data_nxt[0]~40_combout ;
wire \av_ld_byte0_data_nxt[1]~41_combout ;
wire \av_ld_byte0_data_nxt[2]~42_combout ;
wire \av_ld_byte0_data_nxt[3]~43_combout ;
wire \av_ld_byte0_data_nxt[4]~44_combout ;
wire \av_ld_byte0_data_nxt[5]~45_combout ;
wire \av_ld_byte0_data_nxt[6]~46_combout ;
wire \av_ld_byte0_data_nxt[7]~47_combout ;
wire \F_valid~0_combout ;
wire \D_valid~q ;
wire \R_valid~q ;
wire \F_iw[1]~15_combout ;
wire \D_iw[1]~q ;
wire \F_iw[0]~16_combout ;
wire \F_iw[0]~17_combout ;
wire \D_iw[0]~q ;
wire \F_iw[3]~18_combout ;
wire \D_iw[3]~q ;
wire \F_iw[2]~19_combout ;
wire \F_iw[2]~20_combout ;
wire \D_iw[2]~q ;
wire \Equal0~2_combout ;
wire \F_iw[5]~21_combout ;
wire \D_iw[5]~q ;
wire \F_iw[4]~22_combout ;
wire \D_iw[4]~q ;
wire \Equal0~7_combout ;
wire \F_iw[15]~25_combout ;
wire \D_iw[15]~q ;
wire \F_iw[14]~23_combout ;
wire \F_iw[14]~24_combout ;
wire \D_iw[14]~q ;
wire \D_op_opx_rsv63~0_combout ;
wire \F_iw[13]~11_combout ;
wire \D_iw[13]~q ;
wire \F_iw[16]~12_combout ;
wire \D_iw[16]~q ;
wire \F_iw[12]~13_combout ;
wire \F_iw[12]~14_combout ;
wire \D_iw[12]~q ;
wire \Equal62~4_combout ;
wire \Equal62~5_combout ;
wire \Equal62~6_combout ;
wire \D_ctrl_shift_rot~0_combout ;
wire \D_ctrl_shift_logical~0_combout ;
wire \D_ctrl_shift_rot~1_combout ;
wire \Equal62~7_combout ;
wire \D_ctrl_shift_rot~2_combout ;
wire \D_ctrl_shift_rot~3_combout ;
wire \R_ctrl_shift_rot~q ;
wire \E_stall~0_combout ;
wire \E_new_inst~q ;
wire \E_shift_rot_cnt[0]~5_combout ;
wire \D_ctrl_hi_imm16~0_combout ;
wire \D_ctrl_hi_imm16~1_combout ;
wire \R_ctrl_hi_imm16~q ;
wire \D_ctrl_alu_force_xor~14_combout ;
wire \Equal0~17_combout ;
wire \Equal0~11_combout ;
wire \D_ctrl_force_src2_zero~0_combout ;
wire \Equal62~14_combout ;
wire \Equal62~13_combout ;
wire \D_ctrl_force_src2_zero~1_combout ;
wire \Equal62~11_combout ;
wire \D_ctrl_force_src2_zero~2_combout ;
wire \Equal62~9_combout ;
wire \D_ctrl_force_src2_zero~3_combout ;
wire \Equal0~12_combout ;
wire \Equal62~8_combout ;
wire \Equal0~3_combout ;
wire \D_op_cmpge~0_combout ;
wire \D_ctrl_implicit_dst_eretaddr~1_combout ;
wire \Equal62~10_combout ;
wire \D_op_opx_rsv17~0_combout ;
wire \D_ctrl_implicit_dst_eretaddr~2_combout ;
wire \Equal62~2_combout ;
wire \D_op_opx_rsv00~0_combout ;
wire \D_ctrl_implicit_dst_eretaddr~3_combout ;
wire \D_ctrl_implicit_dst_eretaddr~4_combout ;
wire \D_ctrl_implicit_dst_eretaddr~5_combout ;
wire \D_ctrl_implicit_dst_eretaddr~6_combout ;
wire \Equal62~1_combout ;
wire \Equal62~12_combout ;
wire \D_ctrl_implicit_dst_eretaddr~7_combout ;
wire \D_ctrl_implicit_dst_eretaddr~8_combout ;
wire \D_ctrl_implicit_dst_eretaddr~9_combout ;
wire \D_ctrl_implicit_dst_eretaddr~10_combout ;
wire \Equal62~3_combout ;
wire \D_ctrl_implicit_dst_eretaddr~11_combout ;
wire \Equal0~15_combout ;
wire \D_ctrl_implicit_dst_eretaddr~12_combout ;
wire \Equal0~4_combout ;
wire \Equal0~16_combout ;
wire \D_ctrl_force_src2_zero~4_combout ;
wire \D_ctrl_retaddr~0_combout ;
wire \D_ctrl_retaddr~1_combout ;
wire \D_ctrl_retaddr~2_combout ;
wire \D_ctrl_force_src2_zero~5_combout ;
wire \D_ctrl_force_src2_zero~6_combout ;
wire \D_ctrl_force_src2_zero~7_combout ;
wire \D_ctrl_force_src2_zero~8_combout ;
wire \D_ctrl_force_src2_zero~9_combout ;
wire \R_ctrl_force_src2_zero~q ;
wire \R_src2_lo[3]~8_combout ;
wire \F_iw[6]~38_combout ;
wire \F_iw[6]~39_combout ;
wire \D_iw[6]~q ;
wire \D_ctrl_implicit_dst_eretaddr~0_combout ;
wire \D_ctrl_unsigned_lo_imm16~2_combout ;
wire \D_ctrl_unsigned_lo_imm16~5_combout ;
wire \D_ctrl_b_is_dst~0_combout ;
wire \D_ctrl_b_is_dst~1_combout ;
wire \D_ctrl_b_is_dst~2_combout ;
wire \Equal0~13_combout ;
wire \R_src2_use_imm~0_combout ;
wire \R_ctrl_br_nxt~0_combout ;
wire \R_ctrl_br_nxt~1_combout ;
wire \R_src2_use_imm~1_combout ;
wire \R_src2_use_imm~q ;
wire \D_ctrl_src_imm5_shift_rot~0_combout ;
wire \D_ctrl_src_imm5_shift_rot~1_combout ;
wire \R_ctrl_src_imm5_shift_rot~q ;
wire \R_src2_lo~9_combout ;
wire \R_src2_lo[0]~14_combout ;
wire \E_src2[0]~q ;
wire \E_shift_rot_cnt[0]~q ;
wire \E_shift_rot_cnt[0]~6 ;
wire \E_shift_rot_cnt[1]~7_combout ;
wire \F_iw[7]~36_combout ;
wire \F_iw[7]~37_combout ;
wire \D_iw[7]~q ;
wire \R_src2_lo[1]~13_combout ;
wire \E_src2[1]~q ;
wire \E_shift_rot_cnt[1]~q ;
wire \E_shift_rot_cnt[1]~8 ;
wire \E_shift_rot_cnt[2]~9_combout ;
wire \F_iw[8]~34_combout ;
wire \F_iw[8]~35_combout ;
wire \D_iw[8]~q ;
wire \R_src2_lo[2]~12_combout ;
wire \E_src2[2]~q ;
wire \E_shift_rot_cnt[2]~q ;
wire \E_stall~1_combout ;
wire \E_shift_rot_cnt[2]~10 ;
wire \E_shift_rot_cnt[3]~11_combout ;
wire \F_iw[9]~32_combout ;
wire \F_iw[9]~33_combout ;
wire \D_iw[9]~q ;
wire \R_src2_lo[3]~11_combout ;
wire \E_src2[3]~q ;
wire \E_shift_rot_cnt[3]~q ;
wire \E_shift_rot_cnt[3]~12 ;
wire \E_shift_rot_cnt[4]~13_combout ;
wire \F_iw[10]~30_combout ;
wire \F_iw[10]~31_combout ;
wire \D_iw[10]~q ;
wire \R_src2_lo[4]~10_combout ;
wire \E_src2[4]~q ;
wire \E_shift_rot_cnt[4]~q ;
wire \E_stall~2_combout ;
wire \D_ctrl_st~0_combout ;
wire \R_ctrl_st~q ;
wire \D_ctrl_ld_signed~0_combout ;
wire \D_ctrl_ld~2_combout ;
wire \D_ctrl_ld~3_combout ;
wire \R_ctrl_ld~q ;
wire \av_ld_waiting_for_data~q ;
wire \av_ld_waiting_for_data_nxt~0_combout ;
wire \av_ld_waiting_for_data_nxt~1_combout ;
wire \av_ld_aligning_data~q ;
wire \av_ld_align_cycle_nxt[0]~0_combout ;
wire \av_ld_align_cycle[0]~q ;
wire \D_ctrl_mem16~0_combout ;
wire \D_ctrl_mem16~1_combout ;
wire \av_ld_align_cycle_nxt[1]~1_combout ;
wire \av_ld_align_cycle[1]~q ;
wire \av_ld_aligning_data_nxt~0_combout ;
wire \av_ld_aligning_data_nxt~1_combout ;
wire \D_ctrl_mem32~0_combout ;
wire \av_ld_aligning_data_nxt~2_combout ;
wire \E_stall~3_combout ;
wire \E_stall~4_combout ;
wire \E_stall~5_combout ;
wire \E_valid_from_R~0_combout ;
wire \E_valid_from_R~q ;
wire \W_valid~0_combout ;
wire \W_valid~q ;
wire \hbreak_pending_nxt~0_combout ;
wire \hbreak_pending~q ;
wire \wait_for_one_post_bret_inst~0_combout ;
wire \wait_for_one_post_bret_inst~q ;
wire \hbreak_req~0_combout ;
wire \D_ctrl_jmp_direct~0_combout ;
wire \D_ctrl_jmp_direct~1_combout ;
wire \R_ctrl_jmp_direct~q ;
wire \R_ctrl_br~q ;
wire \D_ctrl_retaddr~3_combout ;
wire \D_ctrl_retaddr~4_combout ;
wire \D_ctrl_retaddr~5_combout ;
wire \Equal0~9_combout ;
wire \D_ctrl_retaddr~6_combout ;
wire \D_ctrl_retaddr~7_combout ;
wire \D_ctrl_retaddr~8_combout ;
wire \R_ctrl_retaddr~q ;
wire \R_src1~37_combout ;
wire \R_src1[0]~39_combout ;
wire \E_src1[0]~q ;
wire \D_op_wrctl~combout ;
wire \R_ctrl_wrctl_inst~q ;
wire \E_wrctl_status~0_combout ;
wire \W_estatus_reg_inst_nxt~0_combout ;
wire \W_estatus_reg_inst_nxt~1_combout ;
wire \D_ctrl_exception~3_combout ;
wire \D_ctrl_implicit_dst_eretaddr~16_combout ;
wire \D_ctrl_exception~4_combout ;
wire \D_ctrl_exception~5_combout ;
wire \D_ctrl_implicit_dst_eretaddr~13_combout ;
wire \D_ctrl_exception~0_combout ;
wire \D_ctrl_exception~1_combout ;
wire \D_ctrl_exception~2_combout ;
wire \D_ctrl_exception~6_combout ;
wire \R_ctrl_exception~q ;
wire \W_estatus_reg_inst_nxt~2_combout ;
wire \W_estatus_reg~q ;
wire \W_bstatus_reg_inst_nxt~0_combout ;
wire \W_bstatus_reg_inst_nxt~1_combout ;
wire \D_ctrl_break~0_combout ;
wire \R_ctrl_break~q ;
wire \W_bstatus_reg_inst_nxt~2_combout ;
wire \W_bstatus_reg~q ;
wire \E_wrctl_status~1_combout ;
wire \W_status_reg_pie_inst_nxt~0_combout ;
wire \W_status_reg_pie_inst_nxt~1_combout ;
wire \D_op_eret~combout ;
wire \F_pc_sel_nxt.10~0_combout ;
wire \W_status_reg_pie_inst_nxt~2_combout ;
wire \W_status_reg_pie~q ;
wire \W_ienable_reg_nxt~0_combout ;
wire \W_ienable_reg[0]~0_combout ;
wire \W_ienable_reg[0]~q ;
wire \W_ipending_reg_nxt[0]~0_combout ;
wire \W_ipending_reg[0]~q ;
wire \D_iw[27]~0_combout ;
wire \F_iw[11]~10_combout ;
wire \D_iw[11]~q ;
wire \Equal62~0_combout ;
wire \Equal0~5_combout ;
wire \E_invert_arith_src_msb~0_combout ;
wire \D_ctrl_alu_subtract~2_combout ;
wire \D_ctrl_alu_subtract~3_combout ;
wire \D_ctrl_alu_subtract~4_combout ;
wire \E_alu_sub~0_combout ;
wire \E_alu_sub~q ;
wire \F_iw[18]~26_combout ;
wire \F_iw[18]~27_combout ;
wire \D_iw[18]~q ;
wire \E_src2[7]~15_combout ;
wire \R_src2_lo[12]~0_combout ;
wire \E_src2[12]~q ;
wire \Add1~0_combout ;
wire \R_src1~36_combout ;
wire \E_src1[12]~3_combout ;
wire \F_pc_plus_one[0]~1 ;
wire \F_pc_plus_one[1]~3 ;
wire \F_pc_plus_one[2]~5 ;
wire \F_pc_plus_one[3]~7 ;
wire \F_pc_plus_one[4]~9 ;
wire \F_pc_plus_one[5]~11 ;
wire \F_pc_plus_one[6]~13 ;
wire \F_pc_plus_one[7]~15 ;
wire \F_pc_plus_one[8]~17 ;
wire \F_pc_plus_one[9]~19 ;
wire \F_pc_plus_one[10]~20_combout ;
wire \E_src1[12]~q ;
wire \F_iw[17]~28_combout ;
wire \F_iw[17]~29_combout ;
wire \D_iw[17]~q ;
wire \R_src2_lo[11]~1_combout ;
wire \E_src2[11]~q ;
wire \Add1~1_combout ;
wire \E_src1[11]~4_combout ;
wire \F_pc_plus_one[9]~18_combout ;
wire \E_src1[11]~q ;
wire \R_src2_lo[10]~2_combout ;
wire \E_src2[10]~q ;
wire \Add1~2_combout ;
wire \E_src1[10]~5_combout ;
wire \F_pc_plus_one[8]~16_combout ;
wire \E_src1[10]~q ;
wire \R_src2_lo[9]~3_combout ;
wire \E_src2[9]~q ;
wire \Add1~3_combout ;
wire \E_src1[9]~6_combout ;
wire \F_pc_plus_one[7]~14_combout ;
wire \E_src1[9]~q ;
wire \R_src2_lo[8]~4_combout ;
wire \E_src2[8]~q ;
wire \Add1~4_combout ;
wire \E_src1[8]~7_combout ;
wire \F_pc_plus_one[6]~12_combout ;
wire \E_src1[8]~q ;
wire \R_src2_lo[7]~5_combout ;
wire \E_src2[7]~q ;
wire \Add1~5_combout ;
wire \E_src1[7]~8_combout ;
wire \F_pc_plus_one[5]~10_combout ;
wire \E_src1[7]~q ;
wire \R_src2_lo[6]~6_combout ;
wire \E_src2[6]~q ;
wire \Add1~6_combout ;
wire \E_src1[6]~9_combout ;
wire \F_pc_plus_one[4]~8_combout ;
wire \E_src1[6]~q ;
wire \R_src2_lo[5]~7_combout ;
wire \E_src2[5]~q ;
wire \Add1~7_combout ;
wire \E_src1[5]~10_combout ;
wire \F_pc_plus_one[3]~6_combout ;
wire \E_src1[5]~q ;
wire \Add1~8_combout ;
wire \E_src1[4]~11_combout ;
wire \F_pc_plus_one[2]~4_combout ;
wire \E_src1[4]~q ;
wire \Add1~9_combout ;
wire \E_src1[3]~12_combout ;
wire \F_pc_plus_one[1]~2_combout ;
wire \E_src1[3]~q ;
wire \Add1~10_combout ;
wire \E_src1[2]~13_combout ;
wire \F_pc_plus_one[0]~0_combout ;
wire \E_src1[2]~q ;
wire \Add1~11_combout ;
wire \R_src1[1]~38_combout ;
wire \E_src1[1]~q ;
wire \Add1~12_combout ;
wire \Add1~14_cout ;
wire \Add1~16 ;
wire \Add1~18 ;
wire \Add1~20 ;
wire \Add1~22 ;
wire \Add1~24 ;
wire \Add1~26 ;
wire \Add1~28 ;
wire \Add1~30 ;
wire \Add1~32 ;
wire \Add1~34 ;
wire \Add1~36 ;
wire \Add1~38 ;
wire \Add1~39_combout ;
wire \D_logic_op_raw[1]~0_combout ;
wire \D_ctrl_alu_force_xor~10_combout ;
wire \D_ctrl_alu_force_xor~11_combout ;
wire \D_ctrl_alu_force_xor~13_combout ;
wire \D_ctrl_alu_force_xor~12_combout ;
wire \D_logic_op[1]~0_combout ;
wire \R_logic_op[1]~q ;
wire \D_logic_op[0]~1_combout ;
wire \R_logic_op[0]~q ;
wire \E_logic_result[12]~0_combout ;
wire \Equal0~8_combout ;
wire \Equal0~10_combout ;
wire \D_ctrl_logic~0_combout ;
wire \D_ctrl_logic~combout ;
wire \R_ctrl_logic~q ;
wire \W_alu_result[12]~3_combout ;
wire \D_ctrl_shift_rot_right~0_combout ;
wire \D_ctrl_shift_rot_right~1_combout ;
wire \R_ctrl_shift_rot_right~q ;
wire \E_shift_rot_result_nxt[11]~4_combout ;
wire \E_shift_rot_result[11]~q ;
wire \E_shift_rot_result_nxt[10]~5_combout ;
wire \E_shift_rot_result[10]~q ;
wire \E_shift_rot_result_nxt[9]~6_combout ;
wire \E_shift_rot_result[9]~q ;
wire \E_shift_rot_result_nxt[8]~7_combout ;
wire \E_shift_rot_result[8]~q ;
wire \E_shift_rot_result_nxt[7]~8_combout ;
wire \E_shift_rot_result[7]~q ;
wire \E_shift_rot_result_nxt[6]~9_combout ;
wire \E_shift_rot_result[6]~q ;
wire \E_shift_rot_result_nxt[5]~10_combout ;
wire \E_shift_rot_result[5]~q ;
wire \E_shift_rot_result_nxt[4]~11_combout ;
wire \E_shift_rot_result[4]~q ;
wire \E_shift_rot_result_nxt[3]~12_combout ;
wire \E_shift_rot_result[3]~q ;
wire \E_shift_rot_result_nxt[2]~13_combout ;
wire \E_shift_rot_result[2]~q ;
wire \E_shift_rot_result_nxt[1]~15_combout ;
wire \E_shift_rot_result[1]~q ;
wire \E_shift_rot_result_nxt[0]~16_combout ;
wire \E_shift_rot_result[0]~q ;
wire \R_ctrl_rot_right_nxt~0_combout ;
wire \R_ctrl_rot_right~q ;
wire \D_ctrl_shift_logical~1_combout ;
wire \D_ctrl_shift_logical~2_combout ;
wire \R_ctrl_shift_logical~q ;
wire \E_shift_rot_fill_bit~0_combout ;
wire \E_shift_rot_result_nxt[31]~18_combout ;
wire \R_src1[31]~40_combout ;
wire \E_src1[31]~q ;
wire \E_shift_rot_result[31]~q ;
wire \E_shift_rot_result_nxt[30]~20_combout ;
wire \R_src1[30]~42_combout ;
wire \E_src1[30]~q ;
wire \E_shift_rot_result[30]~q ;
wire \E_shift_rot_result_nxt[29]~22_combout ;
wire \R_src1[29]~43_combout ;
wire \E_src1[29]~q ;
wire \E_shift_rot_result[29]~q ;
wire \E_shift_rot_result_nxt[28]~23_combout ;
wire \R_src1[28]~44_combout ;
wire \E_src1[28]~q ;
wire \E_shift_rot_result[28]~q ;
wire \E_shift_rot_result_nxt[27]~24_combout ;
wire \R_src1[27]~45_combout ;
wire \E_src1[27]~q ;
wire \E_shift_rot_result[27]~q ;
wire \E_shift_rot_result_nxt[26]~25_combout ;
wire \R_src1[26]~46_combout ;
wire \E_src1[26]~q ;
wire \E_shift_rot_result[26]~q ;
wire \E_shift_rot_result_nxt[25]~26_combout ;
wire \R_src1[25]~47_combout ;
wire \E_src1[25]~q ;
wire \E_shift_rot_result[25]~q ;
wire \E_shift_rot_result_nxt[24]~27_combout ;
wire \R_src1[24]~48_combout ;
wire \E_src1[24]~q ;
wire \E_shift_rot_result[24]~q ;
wire \E_shift_rot_result_nxt[23]~28_combout ;
wire \R_src1[23]~49_combout ;
wire \E_src1[23]~q ;
wire \E_shift_rot_result[23]~q ;
wire \E_shift_rot_result_nxt[22]~29_combout ;
wire \R_src1[22]~50_combout ;
wire \E_src1[22]~q ;
wire \E_shift_rot_result[22]~q ;
wire \E_shift_rot_result_nxt[21]~30_combout ;
wire \R_src1[21]~51_combout ;
wire \E_src1[21]~q ;
wire \E_shift_rot_result[21]~q ;
wire \E_shift_rot_result_nxt[20]~31_combout ;
wire \R_src1[20]~52_combout ;
wire \E_src1[20]~q ;
wire \E_shift_rot_result[20]~q ;
wire \E_shift_rot_result_nxt[19]~21_combout ;
wire \R_src1[19]~53_combout ;
wire \E_src1[19]~q ;
wire \E_shift_rot_result[19]~q ;
wire \E_shift_rot_result_nxt[18]~19_combout ;
wire \R_src1[18]~54_combout ;
wire \E_src1[18]~q ;
wire \E_shift_rot_result[18]~q ;
wire \E_shift_rot_result_nxt[17]~17_combout ;
wire \R_src1[17]~55_combout ;
wire \E_src1[17]~q ;
wire \E_shift_rot_result[17]~q ;
wire \E_shift_rot_result_nxt[16]~14_combout ;
wire \R_src1[16]~41_combout ;
wire \E_src1[16]~q ;
wire \E_shift_rot_result[16]~q ;
wire \E_shift_rot_result_nxt[15]~1_combout ;
wire \F_iw[19]~41_combout ;
wire \D_iw[19]~q ;
wire \E_src1[15]~0_combout ;
wire \F_pc_plus_one[10]~21 ;
wire \F_pc_plus_one[11]~23 ;
wire \F_pc_plus_one[12]~25 ;
wire \F_pc_plus_one[13]~26_combout ;
wire \E_src1[15]~q ;
wire \E_shift_rot_result[15]~q ;
wire \E_shift_rot_result_nxt[14]~2_combout ;
wire \E_src1[14]~1_combout ;
wire \F_pc_plus_one[12]~24_combout ;
wire \E_src1[14]~q ;
wire \E_shift_rot_result[14]~q ;
wire \E_shift_rot_result_nxt[13]~3_combout ;
wire \E_src1[13]~2_combout ;
wire \F_pc_plus_one[11]~22_combout ;
wire \E_src1[13]~q ;
wire \E_shift_rot_result[13]~q ;
wire \E_shift_rot_result_nxt[12]~0_combout ;
wire \E_shift_rot_result[12]~q ;
wire \D_op_rdctl~combout ;
wire \R_ctrl_rd_ctl_reg~q ;
wire \Equal0~6_combout ;
wire \D_ctrl_br_cmp~2_combout ;
wire \D_ctrl_br_cmp~5_combout ;
wire \D_ctrl_br_cmp~3_combout ;
wire \D_ctrl_br_cmp~4_combout ;
wire \R_ctrl_br_cmp~q ;
wire \E_alu_result~0_combout ;
wire \F_iw[21]~40_combout ;
wire \D_iw[21]~q ;
wire \R_src2_lo[15]~15_combout ;
wire \E_src2[15]~q ;
wire \Add1~41_combout ;
wire \F_iw[20]~42_combout ;
wire \D_iw[20]~q ;
wire \R_src2_lo[14]~16_combout ;
wire \E_src2[14]~q ;
wire \Add1~42_combout ;
wire \R_src2_lo[13]~17_combout ;
wire \E_src2[13]~q ;
wire \Add1~43_combout ;
wire \Add1~40 ;
wire \Add1~45 ;
wire \Add1~47 ;
wire \Add1~48_combout ;
wire \E_logic_result[15]~1_combout ;
wire \W_alu_result[15]~0_combout ;
wire \Add1~46_combout ;
wire \E_logic_result[14]~2_combout ;
wire \W_alu_result[14]~1_combout ;
wire \Add1~44_combout ;
wire \E_logic_result[13]~3_combout ;
wire \W_alu_result[13]~2_combout ;
wire \Add1~37_combout ;
wire \E_logic_result[11]~4_combout ;
wire \W_alu_result[11]~4_combout ;
wire \Add1~35_combout ;
wire \E_logic_result[10]~5_combout ;
wire \W_alu_result[10]~5_combout ;
wire \Add1~33_combout ;
wire \E_logic_result[9]~6_combout ;
wire \W_alu_result[9]~6_combout ;
wire \Add1~31_combout ;
wire \E_logic_result[8]~7_combout ;
wire \W_alu_result[8]~7_combout ;
wire \Add1~29_combout ;
wire \E_logic_result[7]~8_combout ;
wire \W_alu_result[7]~8_combout ;
wire \Add1~27_combout ;
wire \E_logic_result[6]~9_combout ;
wire \W_alu_result[6]~9_combout ;
wire \Add1~25_combout ;
wire \E_logic_result[5]~10_combout ;
wire \W_alu_result[5]~10_combout ;
wire \Add1~23_combout ;
wire \E_logic_result[4]~11_combout ;
wire \W_alu_result[4]~11_combout ;
wire \Add1~21_combout ;
wire \E_logic_result[3]~12_combout ;
wire \W_alu_result[3]~12_combout ;
wire \Add1~19_combout ;
wire \E_logic_result[2]~13_combout ;
wire \W_alu_result[2]~13_combout ;
wire \d_writedata[24]~0_combout ;
wire \D_ctrl_mem8~0_combout ;
wire \D_ctrl_mem8~1_combout ;
wire \d_writedata[25]~1_combout ;
wire \d_writedata[26]~2_combout ;
wire \d_writedata[27]~3_combout ;
wire \d_writedata[28]~4_combout ;
wire \d_writedata[29]~5_combout ;
wire \d_writedata[30]~6_combout ;
wire \d_writedata[31]~7_combout ;
wire \E_st_stall~combout ;
wire \d_read_nxt~combout ;
wire \D_ctrl_uncond_cti_non_br~0_combout ;
wire \D_ctrl_uncond_cti_non_br~1_combout ;
wire \R_ctrl_uncond_cti_non_br~q ;
wire \Equal0~19_combout ;
wire \R_ctrl_br_uncond~q ;
wire \R_compare_op[1]~q ;
wire \D_logic_op_raw[0]~1_combout ;
wire \R_compare_op[0]~q ;
wire \Equal127~0_combout ;
wire \Equal127~1_combout ;
wire \Equal127~2_combout ;
wire \R_src2_hi[15]~0_combout ;
wire \D_ctrl_unsigned_lo_imm16~3_combout ;
wire \D_ctrl_unsigned_lo_imm16~4_combout ;
wire \R_ctrl_unsigned_lo_imm16~q ;
wire \R_src2_hi[15]~1_combout ;
wire \E_src2[31]~q ;
wire \E_logic_result[31]~14_combout ;
wire \E_logic_result[1]~15_combout ;
wire \Equal127~3_combout ;
wire \Equal127~4_combout ;
wire \E_logic_result[0]~16_combout ;
wire \E_src2[16]~0_combout ;
wire \R_src2_hi~2_combout ;
wire \E_src2[16]~q ;
wire \E_logic_result[16]~17_combout ;
wire \E_src2[30]~1_combout ;
wire \E_src2[30]~q ;
wire \E_logic_result[30]~18_combout ;
wire \E_src2[29]~2_combout ;
wire \E_src2[29]~q ;
wire \E_logic_result[29]~19_combout ;
wire \Equal127~5_combout ;
wire \E_src2[28]~3_combout ;
wire \E_src2[28]~q ;
wire \E_logic_result[28]~20_combout ;
wire \E_src2[27]~4_combout ;
wire \E_src2[27]~q ;
wire \E_logic_result[27]~21_combout ;
wire \E_src2[26]~5_combout ;
wire \E_src2[26]~q ;
wire \E_logic_result[26]~22_combout ;
wire \E_src2[25]~6_combout ;
wire \E_src2[25]~q ;
wire \E_logic_result[25]~23_combout ;
wire \Equal127~6_combout ;
wire \E_src2[24]~7_combout ;
wire \E_src2[24]~q ;
wire \E_logic_result[24]~24_combout ;
wire \E_src2[23]~8_combout ;
wire \E_src2[23]~q ;
wire \E_logic_result[23]~25_combout ;
wire \E_src2[22]~9_combout ;
wire \E_src2[22]~q ;
wire \E_logic_result[22]~26_combout ;
wire \E_src2[21]~10_combout ;
wire \E_src2[21]~q ;
wire \E_logic_result[21]~27_combout ;
wire \Equal127~7_combout ;
wire \E_src2[20]~11_combout ;
wire \E_src2[20]~q ;
wire \E_logic_result[20]~28_combout ;
wire \E_src2[19]~12_combout ;
wire \E_src2[19]~q ;
wire \E_logic_result[19]~29_combout ;
wire \E_src2[18]~13_combout ;
wire \E_src2[18]~q ;
wire \E_logic_result[18]~30_combout ;
wire \E_src2[17]~14_combout ;
wire \E_src2[17]~q ;
wire \E_logic_result[17]~31_combout ;
wire \Equal127~8_combout ;
wire \Equal127~9_combout ;
wire \E_cmp_result~0_combout ;
wire \E_invert_arith_src_msb~1_combout ;
wire \E_invert_arith_src_msb~2_combout ;
wire \E_invert_arith_src_msb~q ;
wire \Add1~50_combout ;
wire \E_arith_src1[31]~combout ;
wire \Add1~51_combout ;
wire \Add1~52_combout ;
wire \Add1~53_combout ;
wire \Add1~54_combout ;
wire \Add1~55_combout ;
wire \Add1~56_combout ;
wire \Add1~57_combout ;
wire \Add1~58_combout ;
wire \Add1~59_combout ;
wire \Add1~60_combout ;
wire \Add1~61_combout ;
wire \Add1~62_combout ;
wire \Add1~63_combout ;
wire \Add1~64_combout ;
wire \Add1~65_combout ;
wire \Add1~49 ;
wire \Add1~67 ;
wire \Add1~69 ;
wire \Add1~71 ;
wire \Add1~73 ;
wire \Add1~75 ;
wire \Add1~77 ;
wire \Add1~79 ;
wire \Add1~81 ;
wire \Add1~83 ;
wire \Add1~85 ;
wire \Add1~87 ;
wire \Add1~89 ;
wire \Add1~91 ;
wire \Add1~93 ;
wire \Add1~95 ;
wire \Add1~97 ;
wire \Add1~98_combout ;
wire \E_cmp_result~1_combout ;
wire \W_cmp_result~q ;
wire \F_pc_sel_nxt~0_combout ;
wire \F_pc_no_crst_nxt[10]~0_combout ;
wire \F_pc_no_crst_nxt[9]~1_combout ;
wire \F_pc_no_crst_nxt[9]~2_combout ;
wire \F_pc_no_crst_nxt[8]~3_combout ;
wire \F_pc_no_crst_nxt[7]~4_combout ;
wire \F_pc_no_crst_nxt[6]~5_combout ;
wire \F_pc_no_crst_nxt[5]~6_combout ;
wire \F_pc_no_crst_nxt[4]~7_combout ;
wire \F_pc_no_crst_nxt[3]~8_combout ;
wire \F_pc_no_crst_nxt[2]~9_combout ;
wire \F_pc_no_crst_nxt[1]~10_combout ;
wire \F_pc_no_crst_nxt[0]~11_combout ;
wire \F_pc_no_crst_nxt[13]~12_combout ;
wire \F_pc_no_crst_nxt[13]~13_combout ;
wire \F_pc_no_crst_nxt[12]~14_combout ;
wire \F_pc_no_crst_nxt[11]~15_combout ;
wire \i_read_nxt~0_combout ;
wire \hbreak_enabled~0_combout ;
wire \Add1~15_combout ;
wire \Add1~17_combout ;
wire \E_mem_byte_en[0]~0_combout ;
wire \d_byteenable[3]~0_combout ;
wire \E_st_data[22]~0_combout ;
wire \E_mem_byte_en[2]~1_combout ;
wire \E_st_data[23]~1_combout ;
wire \E_mem_byte_en[3]~2_combout ;
wire \E_st_data[11]~2_combout ;
wire \E_mem_byte_en[1]~3_combout ;
wire \E_st_data[13]~3_combout ;
wire \E_st_data[16]~4_combout ;
wire \E_st_data[12]~5_combout ;
wire \E_st_data[14]~6_combout ;
wire \E_st_data[15]~7_combout ;
wire \E_st_data[18]~8_combout ;
wire \E_st_data[17]~9_combout ;
wire \E_st_data[10]~10_combout ;
wire \E_st_data[9]~11_combout ;
wire \E_st_data[8]~12_combout ;
wire \E_st_data[21]~13_combout ;
wire \E_st_data[19]~14_combout ;
wire \E_st_data[20]~15_combout ;


nios_mcu_nios_mcu_nios_cpu_cpu_nios2_oci the_nios_mcu_nios_cpu_cpu_nios2_oci(
	.sr_0(sr_0),
	.jtag_break(\the_nios_mcu_nios_cpu_cpu_nios2_oci|the_nios_mcu_nios_cpu_cpu_nios2_oci_debug|jtag_break~q ),
	.readdata_0(readdata_0),
	.readdata_1(readdata_1),
	.readdata_3(readdata_3),
	.readdata_2(readdata_2),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.r_sync_rst(r_sync_rst),
	.m0_write(m0_write),
	.saved_grant_0(saved_grant_0),
	.waitrequest(debug_mem_slave_waitrequest),
	.mem_used_1(mem_used_1),
	.WideOr1(WideOr12),
	.rf_source_valid(rf_source_valid),
	.hbreak_enabled(hbreak_enabled1),
	.address_nxt({src_data_46,src_data_45,src_data_44,src_data_43,src_data_42,src_data_41,src_data_40,src_data_39,src_data_38}),
	.r_early_rst(r_early_rst),
	.oci_ienable_0(\the_nios_mcu_nios_cpu_cpu_nios2_oci|the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_ienable[0]~q ),
	.oci_single_step_mode(\the_nios_mcu_nios_cpu_cpu_nios2_oci|the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_single_step_mode~q ),
	.readdata_22(readdata_22),
	.readdata_23(readdata_23),
	.readdata_24(readdata_24),
	.readdata_25(readdata_25),
	.readdata_26(readdata_26),
	.readdata_11(readdata_11),
	.readdata_13(readdata_13),
	.readdata_16(readdata_16),
	.readdata_12(readdata_12),
	.readdata_5(readdata_5),
	.readdata_4(readdata_4),
	.readdata_14(readdata_14),
	.readdata_15(readdata_15),
	.readdata_18(readdata_18),
	.readdata_17(readdata_17),
	.readdata_10(readdata_10),
	.readdata_9(readdata_9),
	.readdata_8(readdata_8),
	.readdata_7(readdata_7),
	.readdata_6(readdata_6),
	.readdata_21(readdata_21),
	.readdata_19(readdata_19),
	.readdata_20(readdata_20),
	.debugaccess_nxt(src_payload11),
	.writedata_nxt({src_payload43,src_payload42,src_payload41,src_payload40,src_payload39,src_payload20,src_payload19,src_payload18,src_payload17,src_payload16,src_payload36,src_payload38,src_payload37,src_payload29,src_payload30,src_payload23,src_payload28,src_payload27,src_payload22,
src_payload24,src_payload21,src_payload31,src_payload32,src_payload33,src_payload34,src_payload35,src_payload25,src_payload26,src_payload14,src_payload15,src_payload13,src_payload12}),
	.byteenable_nxt({src_data_35,src_data_34,src_data_33,src_data_32}),
	.readdata_27(readdata_27),
	.readdata_28(readdata_28),
	.readdata_29(readdata_29),
	.readdata_30(readdata_30),
	.readdata_31(readdata_31),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_1(state_1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3),
	.irf_reg_0_2(irf_reg_0_2),
	.irf_reg_1_2(irf_reg_1_2),
	.clk_clk(clk_clk));

nios_mcu_nios_mcu_nios_cpu_cpu_register_bank_b_module nios_mcu_nios_cpu_cpu_register_bank_b(
	.q_b_0(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.q_b_1(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_2(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.q_b_3(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.q_b_4(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.q_b_5(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.q_b_6(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.q_b_7(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.q_b_12(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ),
	.q_b_11(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ),
	.q_b_10(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ),
	.q_b_9(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ),
	.q_b_8(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ),
	.q_b_15(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ),
	.q_b_14(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ),
	.q_b_13(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ),
	.q_b_31(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[31] ),
	.q_b_16(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[16] ),
	.q_b_30(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[30] ),
	.q_b_29(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[29] ),
	.q_b_28(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[28] ),
	.q_b_27(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[27] ),
	.q_b_26(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[26] ),
	.q_b_25(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[25] ),
	.q_b_24(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[24] ),
	.q_b_23(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[23] ),
	.q_b_22(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[22] ),
	.q_b_21(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[21] ),
	.q_b_20(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[20] ),
	.q_b_19(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[19] ),
	.q_b_18(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[18] ),
	.q_b_17(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[17] ),
	.W_rf_wren(\W_rf_wren~combout ),
	.W_rf_wr_data_0(\W_rf_wr_data[0]~2_combout ),
	.R_dst_regnum_0(\R_dst_regnum[0]~q ),
	.R_dst_regnum_1(\R_dst_regnum[1]~q ),
	.R_dst_regnum_2(\R_dst_regnum[2]~q ),
	.R_dst_regnum_3(\R_dst_regnum[3]~q ),
	.R_dst_regnum_4(\R_dst_regnum[4]~q ),
	.D_iw_22(\D_iw[22]~q ),
	.D_iw_23(\D_iw[23]~q ),
	.D_iw_24(\D_iw[24]~q ),
	.D_iw_25(\D_iw[25]~q ),
	.D_iw_26(\D_iw[26]~q ),
	.W_rf_wr_data_1(\W_rf_wr_data[1]~3_combout ),
	.W_rf_wr_data_2(\W_rf_wr_data[2]~4_combout ),
	.W_rf_wr_data_3(\W_rf_wr_data[3]~5_combout ),
	.W_rf_wr_data_4(\W_rf_wr_data[4]~6_combout ),
	.W_rf_wr_data_5(\W_rf_wr_data[5]~7_combout ),
	.W_rf_wr_data_6(\W_rf_wr_data[6]~8_combout ),
	.W_rf_wr_data_7(\W_rf_wr_data[7]~9_combout ),
	.W_rf_wr_data_12(\W_rf_wr_data[12]~10_combout ),
	.W_rf_wr_data_11(\W_rf_wr_data[11]~11_combout ),
	.W_rf_wr_data_10(\W_rf_wr_data[10]~12_combout ),
	.W_rf_wr_data_9(\W_rf_wr_data[9]~13_combout ),
	.W_rf_wr_data_8(\W_rf_wr_data[8]~14_combout ),
	.W_rf_wr_data_15(\W_rf_wr_data[15]~15_combout ),
	.W_rf_wr_data_14(\W_rf_wr_data[14]~16_combout ),
	.W_rf_wr_data_13(\W_rf_wr_data[13]~17_combout ),
	.W_rf_wr_data_31(\W_rf_wr_data[31]~18_combout ),
	.W_rf_wr_data_16(\W_rf_wr_data[16]~19_combout ),
	.W_rf_wr_data_30(\W_rf_wr_data[30]~20_combout ),
	.W_rf_wr_data_29(\W_rf_wr_data[29]~21_combout ),
	.W_rf_wr_data_28(\W_rf_wr_data[28]~22_combout ),
	.W_rf_wr_data_27(\W_rf_wr_data[27]~23_combout ),
	.W_rf_wr_data_26(\W_rf_wr_data[26]~24_combout ),
	.W_rf_wr_data_25(\W_rf_wr_data[25]~25_combout ),
	.W_rf_wr_data_24(\W_rf_wr_data[24]~26_combout ),
	.W_rf_wr_data_23(\W_rf_wr_data[23]~27_combout ),
	.W_rf_wr_data_22(\W_rf_wr_data[22]~28_combout ),
	.W_rf_wr_data_21(\W_rf_wr_data[21]~29_combout ),
	.W_rf_wr_data_20(\W_rf_wr_data[20]~30_combout ),
	.W_rf_wr_data_19(\W_rf_wr_data[19]~31_combout ),
	.W_rf_wr_data_18(\W_rf_wr_data[18]~32_combout ),
	.W_rf_wr_data_17(\W_rf_wr_data[17]~33_combout ),
	.clk_clk(clk_clk));

nios_mcu_nios_mcu_nios_cpu_cpu_register_bank_a_module nios_mcu_nios_cpu_cpu_register_bank_a(
	.q_b_12(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[12] ),
	.q_b_11(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[11] ),
	.q_b_10(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[10] ),
	.q_b_9(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[9] ),
	.q_b_8(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[8] ),
	.q_b_7(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[7] ),
	.q_b_6(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[6] ),
	.q_b_5(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[5] ),
	.q_b_4(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[4] ),
	.q_b_3(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[3] ),
	.q_b_2(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[2] ),
	.q_b_1(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_0(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[0] ),
	.q_b_15(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[15] ),
	.q_b_14(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[14] ),
	.q_b_13(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[13] ),
	.q_b_31(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[31] ),
	.q_b_16(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[16] ),
	.q_b_30(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[30] ),
	.q_b_29(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[29] ),
	.q_b_28(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[28] ),
	.q_b_27(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[27] ),
	.q_b_26(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[26] ),
	.q_b_25(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[25] ),
	.q_b_24(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[24] ),
	.q_b_23(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[23] ),
	.q_b_22(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[22] ),
	.q_b_21(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[21] ),
	.q_b_20(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[20] ),
	.q_b_19(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[19] ),
	.q_b_18(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[18] ),
	.q_b_17(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[17] ),
	.W_rf_wren(\W_rf_wren~combout ),
	.W_rf_wr_data_0(\W_rf_wr_data[0]~2_combout ),
	.R_dst_regnum_0(\R_dst_regnum[0]~q ),
	.R_dst_regnum_1(\R_dst_regnum[1]~q ),
	.R_dst_regnum_2(\R_dst_regnum[2]~q ),
	.R_dst_regnum_3(\R_dst_regnum[3]~q ),
	.R_dst_regnum_4(\R_dst_regnum[4]~q ),
	.W_rf_wr_data_1(\W_rf_wr_data[1]~3_combout ),
	.W_rf_wr_data_2(\W_rf_wr_data[2]~4_combout ),
	.W_rf_wr_data_3(\W_rf_wr_data[3]~5_combout ),
	.W_rf_wr_data_4(\W_rf_wr_data[4]~6_combout ),
	.W_rf_wr_data_5(\W_rf_wr_data[5]~7_combout ),
	.W_rf_wr_data_6(\W_rf_wr_data[6]~8_combout ),
	.W_rf_wr_data_7(\W_rf_wr_data[7]~9_combout ),
	.W_rf_wr_data_12(\W_rf_wr_data[12]~10_combout ),
	.D_iw_27(\D_iw[27]~q ),
	.D_iw_28(\D_iw[28]~q ),
	.D_iw_29(\D_iw[29]~q ),
	.D_iw_30(\D_iw[30]~q ),
	.D_iw_31(\D_iw[31]~q ),
	.W_rf_wr_data_11(\W_rf_wr_data[11]~11_combout ),
	.W_rf_wr_data_10(\W_rf_wr_data[10]~12_combout ),
	.W_rf_wr_data_9(\W_rf_wr_data[9]~13_combout ),
	.W_rf_wr_data_8(\W_rf_wr_data[8]~14_combout ),
	.W_rf_wr_data_15(\W_rf_wr_data[15]~15_combout ),
	.W_rf_wr_data_14(\W_rf_wr_data[14]~16_combout ),
	.W_rf_wr_data_13(\W_rf_wr_data[13]~17_combout ),
	.W_rf_wr_data_31(\W_rf_wr_data[31]~18_combout ),
	.W_rf_wr_data_16(\W_rf_wr_data[16]~19_combout ),
	.W_rf_wr_data_30(\W_rf_wr_data[30]~20_combout ),
	.W_rf_wr_data_29(\W_rf_wr_data[29]~21_combout ),
	.W_rf_wr_data_28(\W_rf_wr_data[28]~22_combout ),
	.W_rf_wr_data_27(\W_rf_wr_data[27]~23_combout ),
	.W_rf_wr_data_26(\W_rf_wr_data[26]~24_combout ),
	.W_rf_wr_data_25(\W_rf_wr_data[25]~25_combout ),
	.W_rf_wr_data_24(\W_rf_wr_data[24]~26_combout ),
	.W_rf_wr_data_23(\W_rf_wr_data[23]~27_combout ),
	.W_rf_wr_data_22(\W_rf_wr_data[22]~28_combout ),
	.W_rf_wr_data_21(\W_rf_wr_data[21]~29_combout ),
	.W_rf_wr_data_20(\W_rf_wr_data[20]~30_combout ),
	.W_rf_wr_data_19(\W_rf_wr_data[19]~31_combout ),
	.W_rf_wr_data_18(\W_rf_wr_data[18]~32_combout ),
	.W_rf_wr_data_17(\W_rf_wr_data[17]~33_combout ),
	.clk_clk(clk_clk));

dffeas \W_alu_result[0] (
	.clk(clk_clk),
	.d(\W_alu_result[0]~14_combout ),
	.asdata(\E_shift_rot_result[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[0]~q ),
	.prn(vcc));
defparam \W_alu_result[0] .is_wysiwyg = "true";
defparam \W_alu_result[0] .power_up = "low";

dffeas \W_alu_result[1] (
	.clk(clk_clk),
	.d(\W_alu_result[1]~15_combout ),
	.asdata(\E_shift_rot_result[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[1]~q ),
	.prn(vcc));
defparam \W_alu_result[1] .is_wysiwyg = "true";
defparam \W_alu_result[1] .power_up = "low";

dffeas \av_ld_byte1_data[0] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[0]~0_combout ),
	.asdata(\av_ld_byte2_data[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[0]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[0] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[0] .power_up = "low";

cycloneive_lcell_comb \Add1~66 (
	.dataa(\Add1~65_combout ),
	.datab(\E_src1[16]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~49 ),
	.combout(\Add1~66_combout ),
	.cout(\Add1~67 ));
defparam \Add1~66 .lut_mask = 16'h967F;
defparam \Add1~66 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~68 (
	.dataa(\Add1~64_combout ),
	.datab(\E_src1[17]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~67 ),
	.combout(\Add1~68_combout ),
	.cout(\Add1~69 ));
defparam \Add1~68 .lut_mask = 16'h96EF;
defparam \Add1~68 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~70 (
	.dataa(\Add1~63_combout ),
	.datab(\E_src1[18]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~69 ),
	.combout(\Add1~70_combout ),
	.cout(\Add1~71 ));
defparam \Add1~70 .lut_mask = 16'h967F;
defparam \Add1~70 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~72 (
	.dataa(\Add1~62_combout ),
	.datab(\E_src1[19]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~71 ),
	.combout(\Add1~72_combout ),
	.cout(\Add1~73 ));
defparam \Add1~72 .lut_mask = 16'h96EF;
defparam \Add1~72 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~74 (
	.dataa(\Add1~61_combout ),
	.datab(\E_src1[20]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~73 ),
	.combout(\Add1~74_combout ),
	.cout(\Add1~75 ));
defparam \Add1~74 .lut_mask = 16'h967F;
defparam \Add1~74 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~76 (
	.dataa(\Add1~60_combout ),
	.datab(\E_src1[21]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~75 ),
	.combout(\Add1~76_combout ),
	.cout(\Add1~77 ));
defparam \Add1~76 .lut_mask = 16'h96EF;
defparam \Add1~76 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~78 (
	.dataa(\Add1~59_combout ),
	.datab(\E_src1[22]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~77 ),
	.combout(\Add1~78_combout ),
	.cout(\Add1~79 ));
defparam \Add1~78 .lut_mask = 16'h967F;
defparam \Add1~78 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~80 (
	.dataa(\Add1~58_combout ),
	.datab(\E_src1[23]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~79 ),
	.combout(\Add1~80_combout ),
	.cout(\Add1~81 ));
defparam \Add1~80 .lut_mask = 16'h96EF;
defparam \Add1~80 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~82 (
	.dataa(\Add1~57_combout ),
	.datab(\E_src1[24]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~81 ),
	.combout(\Add1~82_combout ),
	.cout(\Add1~83 ));
defparam \Add1~82 .lut_mask = 16'h967F;
defparam \Add1~82 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~84 (
	.dataa(\Add1~56_combout ),
	.datab(\E_src1[25]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~83 ),
	.combout(\Add1~84_combout ),
	.cout(\Add1~85 ));
defparam \Add1~84 .lut_mask = 16'h96EF;
defparam \Add1~84 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~86 (
	.dataa(\Add1~55_combout ),
	.datab(\E_src1[26]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~85 ),
	.combout(\Add1~86_combout ),
	.cout(\Add1~87 ));
defparam \Add1~86 .lut_mask = 16'h967F;
defparam \Add1~86 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~88 (
	.dataa(\Add1~54_combout ),
	.datab(\E_src1[27]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~87 ),
	.combout(\Add1~88_combout ),
	.cout(\Add1~89 ));
defparam \Add1~88 .lut_mask = 16'h96EF;
defparam \Add1~88 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~90 (
	.dataa(\Add1~53_combout ),
	.datab(\E_src1[28]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~89 ),
	.combout(\Add1~90_combout ),
	.cout(\Add1~91 ));
defparam \Add1~90 .lut_mask = 16'h967F;
defparam \Add1~90 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~92 (
	.dataa(\Add1~52_combout ),
	.datab(\E_src1[29]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~91 ),
	.combout(\Add1~92_combout ),
	.cout(\Add1~93 ));
defparam \Add1~92 .lut_mask = 16'h96EF;
defparam \Add1~92 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~94 (
	.dataa(\Add1~51_combout ),
	.datab(\E_src1[30]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~93 ),
	.combout(\Add1~94_combout ),
	.cout(\Add1~95 ));
defparam \Add1~94 .lut_mask = 16'h967F;
defparam \Add1~94 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~96 (
	.dataa(\Add1~50_combout ),
	.datab(\E_arith_src1[31]~combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~95 ),
	.combout(\Add1~96_combout ),
	.cout(\Add1~97 ));
defparam \Add1~96 .lut_mask = 16'h96EF;
defparam \Add1~96 .sum_lutc_input = "cin";

cycloneive_lcell_comb \W_alu_result[0]~14 (
	.dataa(\Add1~15_combout ),
	.datab(\E_logic_result[0]~16_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[0]~14_combout ),
	.cout());
defparam \W_alu_result[0]~14 .lut_mask = 16'hAACC;
defparam \W_alu_result[0]~14 .sum_lutc_input = "datac";

dffeas \av_ld_byte1_data[4] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[4]~4_combout ),
	.asdata(\av_ld_byte2_data[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[4]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[4] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[4] .power_up = "low";

dffeas \av_ld_byte1_data[3] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[3]~5_combout ),
	.asdata(\av_ld_byte2_data[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[3]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[3] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[3] .power_up = "low";

dffeas \av_ld_byte1_data[2] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[2]~6_combout ),
	.asdata(\av_ld_byte2_data[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[2]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[2] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[2] .power_up = "low";

dffeas \av_ld_byte1_data[1] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[1]~7_combout ),
	.asdata(\av_ld_byte2_data[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[1]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[1] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[1] .power_up = "low";

dffeas \av_ld_byte1_data[7] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[7]~1_combout ),
	.asdata(\av_ld_byte2_data[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[7]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[7] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[7] .power_up = "low";

dffeas \av_ld_byte1_data[6] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[6]~2_combout ),
	.asdata(\av_ld_byte2_data[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[6]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[6] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[6] .power_up = "low";

dffeas \av_ld_byte1_data[5] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[5]~3_combout ),
	.asdata(\av_ld_byte2_data[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(\av_ld_byte1_data_en~0_combout ),
	.q(\av_ld_byte1_data[5]~q ),
	.prn(vcc));
defparam \av_ld_byte1_data[5] .is_wysiwyg = "true";
defparam \av_ld_byte1_data[5] .power_up = "low";

cycloneive_lcell_comb \W_alu_result[1]~15 (
	.dataa(\Add1~17_combout ),
	.datab(\E_logic_result[1]~15_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[1]~15_combout ),
	.cout());
defparam \W_alu_result[1]~15 .lut_mask = 16'hAACC;
defparam \W_alu_result[1]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte1_data[0]~0 (
	.dataa(src_data_8),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[0]~0_combout ),
	.cout());
defparam \av_ld_byte1_data[0]~0 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[0]~0 .sum_lutc_input = "datac";

dffeas \av_ld_byte2_data[0] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data[0]~0_combout ),
	.asdata(\av_ld_byte3_data[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[0]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[0] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[0] .power_up = "low";

cycloneive_lcell_comb \av_ld_byte1_data[4]~4 (
	.dataa(src_data_12),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[4]~4_combout ),
	.cout());
defparam \av_ld_byte1_data[4]~4 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[4]~4 .sum_lutc_input = "datac";

dffeas \av_ld_byte2_data[4] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data[4]~4_combout ),
	.asdata(\av_ld_byte3_data[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[4]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[4] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[4] .power_up = "low";

cycloneive_lcell_comb \av_ld_byte1_data[3]~5 (
	.dataa(src_data_11),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[3]~5_combout ),
	.cout());
defparam \av_ld_byte1_data[3]~5 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[3]~5 .sum_lutc_input = "datac";

dffeas \av_ld_byte2_data[3] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data[3]~5_combout ),
	.asdata(\av_ld_byte3_data[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[3]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[3] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[3] .power_up = "low";

cycloneive_lcell_comb \av_ld_byte1_data[2]~6 (
	.dataa(src_data_10),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[2]~6_combout ),
	.cout());
defparam \av_ld_byte1_data[2]~6 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[2]~6 .sum_lutc_input = "datac";

dffeas \av_ld_byte2_data[2] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data[2]~6_combout ),
	.asdata(\av_ld_byte3_data[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[2]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[2] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[2] .power_up = "low";

cycloneive_lcell_comb \av_ld_byte1_data[1]~7 (
	.dataa(src_data_9),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[1]~7_combout ),
	.cout());
defparam \av_ld_byte1_data[1]~7 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[1]~7 .sum_lutc_input = "datac";

dffeas \av_ld_byte2_data[1] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data[1]~7_combout ),
	.asdata(\av_ld_byte3_data[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[1]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[1] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[1] .power_up = "low";

cycloneive_lcell_comb \av_ld_byte1_data[7]~1 (
	.dataa(src_data_15),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[7]~1_combout ),
	.cout());
defparam \av_ld_byte1_data[7]~1 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[7]~1 .sum_lutc_input = "datac";

dffeas \av_ld_byte2_data[7] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data[7]~1_combout ),
	.asdata(\av_ld_byte3_data[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[7]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[7] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[7] .power_up = "low";

cycloneive_lcell_comb \av_ld_byte1_data[6]~2 (
	.dataa(src_data_14),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[6]~2_combout ),
	.cout());
defparam \av_ld_byte1_data[6]~2 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[6]~2 .sum_lutc_input = "datac";

dffeas \av_ld_byte2_data[6] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data[6]~2_combout ),
	.asdata(\av_ld_byte3_data[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[6]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[6] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[6] .power_up = "low";

cycloneive_lcell_comb \av_ld_byte1_data[5]~3 (
	.dataa(src_data_13),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte1_data[5]~3_combout ),
	.cout());
defparam \av_ld_byte1_data[5]~3 .lut_mask = 16'hAACC;
defparam \av_ld_byte1_data[5]~3 .sum_lutc_input = "datac";

dffeas \av_ld_byte2_data[5] (
	.clk(clk_clk),
	.d(\av_ld_byte2_data[5]~3_combout ),
	.asdata(\av_ld_byte3_data[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\av_ld_rshift8~1_combout ),
	.ena(vcc),
	.q(\av_ld_byte2_data[5]~q ),
	.prn(vcc));
defparam \av_ld_byte2_data[5] .is_wysiwyg = "true";
defparam \av_ld_byte2_data[5] .power_up = "low";

cycloneive_lcell_comb \av_ld_byte2_data[0]~0 (
	.dataa(src_data_16),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[0]~0_combout ),
	.cout());
defparam \av_ld_byte2_data[0]~0 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[0]~0 .sum_lutc_input = "datac";

dffeas \W_alu_result[31] (
	.clk(clk_clk),
	.d(\W_alu_result[31]~16_combout ),
	.asdata(\E_shift_rot_result[31]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[31]~q ),
	.prn(vcc));
defparam \W_alu_result[31] .is_wysiwyg = "true";
defparam \W_alu_result[31] .power_up = "low";

dffeas \W_alu_result[16] (
	.clk(clk_clk),
	.d(\W_alu_result[16]~17_combout ),
	.asdata(\E_shift_rot_result[16]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[16]~q ),
	.prn(vcc));
defparam \W_alu_result[16] .is_wysiwyg = "true";
defparam \W_alu_result[16] .power_up = "low";

dffeas \W_alu_result[30] (
	.clk(clk_clk),
	.d(\W_alu_result[30]~18_combout ),
	.asdata(\E_shift_rot_result[30]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[30]~q ),
	.prn(vcc));
defparam \W_alu_result[30] .is_wysiwyg = "true";
defparam \W_alu_result[30] .power_up = "low";

dffeas \W_alu_result[29] (
	.clk(clk_clk),
	.d(\W_alu_result[29]~19_combout ),
	.asdata(\E_shift_rot_result[29]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[29]~q ),
	.prn(vcc));
defparam \W_alu_result[29] .is_wysiwyg = "true";
defparam \W_alu_result[29] .power_up = "low";

dffeas \W_alu_result[28] (
	.clk(clk_clk),
	.d(\W_alu_result[28]~20_combout ),
	.asdata(\E_shift_rot_result[28]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[28]~q ),
	.prn(vcc));
defparam \W_alu_result[28] .is_wysiwyg = "true";
defparam \W_alu_result[28] .power_up = "low";

dffeas \W_alu_result[27] (
	.clk(clk_clk),
	.d(\W_alu_result[27]~21_combout ),
	.asdata(\E_shift_rot_result[27]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[27]~q ),
	.prn(vcc));
defparam \W_alu_result[27] .is_wysiwyg = "true";
defparam \W_alu_result[27] .power_up = "low";

dffeas \W_alu_result[26] (
	.clk(clk_clk),
	.d(\W_alu_result[26]~22_combout ),
	.asdata(\E_shift_rot_result[26]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[26]~q ),
	.prn(vcc));
defparam \W_alu_result[26] .is_wysiwyg = "true";
defparam \W_alu_result[26] .power_up = "low";

dffeas \W_alu_result[25] (
	.clk(clk_clk),
	.d(\W_alu_result[25]~23_combout ),
	.asdata(\E_shift_rot_result[25]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[25]~q ),
	.prn(vcc));
defparam \W_alu_result[25] .is_wysiwyg = "true";
defparam \W_alu_result[25] .power_up = "low";

dffeas \W_alu_result[24] (
	.clk(clk_clk),
	.d(\W_alu_result[24]~24_combout ),
	.asdata(\E_shift_rot_result[24]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[24]~q ),
	.prn(vcc));
defparam \W_alu_result[24] .is_wysiwyg = "true";
defparam \W_alu_result[24] .power_up = "low";

dffeas \W_alu_result[23] (
	.clk(clk_clk),
	.d(\W_alu_result[23]~25_combout ),
	.asdata(\E_shift_rot_result[23]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[23]~q ),
	.prn(vcc));
defparam \W_alu_result[23] .is_wysiwyg = "true";
defparam \W_alu_result[23] .power_up = "low";

dffeas \W_alu_result[22] (
	.clk(clk_clk),
	.d(\W_alu_result[22]~26_combout ),
	.asdata(\E_shift_rot_result[22]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[22]~q ),
	.prn(vcc));
defparam \W_alu_result[22] .is_wysiwyg = "true";
defparam \W_alu_result[22] .power_up = "low";

dffeas \W_alu_result[21] (
	.clk(clk_clk),
	.d(\W_alu_result[21]~27_combout ),
	.asdata(\E_shift_rot_result[21]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[21]~q ),
	.prn(vcc));
defparam \W_alu_result[21] .is_wysiwyg = "true";
defparam \W_alu_result[21] .power_up = "low";

dffeas \W_alu_result[20] (
	.clk(clk_clk),
	.d(\W_alu_result[20]~28_combout ),
	.asdata(\E_shift_rot_result[20]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[20]~q ),
	.prn(vcc));
defparam \W_alu_result[20] .is_wysiwyg = "true";
defparam \W_alu_result[20] .power_up = "low";

dffeas \W_alu_result[19] (
	.clk(clk_clk),
	.d(\W_alu_result[19]~29_combout ),
	.asdata(\E_shift_rot_result[19]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[19]~q ),
	.prn(vcc));
defparam \W_alu_result[19] .is_wysiwyg = "true";
defparam \W_alu_result[19] .power_up = "low";

dffeas \W_alu_result[18] (
	.clk(clk_clk),
	.d(\W_alu_result[18]~30_combout ),
	.asdata(\E_shift_rot_result[18]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[18]~q ),
	.prn(vcc));
defparam \W_alu_result[18] .is_wysiwyg = "true";
defparam \W_alu_result[18] .power_up = "low";

dffeas \W_alu_result[17] (
	.clk(clk_clk),
	.d(\W_alu_result[17]~31_combout ),
	.asdata(\E_shift_rot_result[17]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(\W_alu_result[17]~q ),
	.prn(vcc));
defparam \W_alu_result[17] .is_wysiwyg = "true";
defparam \W_alu_result[17] .power_up = "low";

cycloneive_lcell_comb \av_ld_byte2_data[4]~4 (
	.dataa(src_data_20),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[4]~4_combout ),
	.cout());
defparam \av_ld_byte2_data[4]~4 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte2_data[3]~5 (
	.dataa(src_data_19),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[3]~5_combout ),
	.cout());
defparam \av_ld_byte2_data[3]~5 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[3]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte2_data[2]~6 (
	.dataa(src_data_18),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[2]~6_combout ),
	.cout());
defparam \av_ld_byte2_data[2]~6 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[2]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte2_data[1]~7 (
	.dataa(src_data_17),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[1]~7_combout ),
	.cout());
defparam \av_ld_byte2_data[1]~7 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[1]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte2_data[7]~1 (
	.dataa(src_data_23),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[7]~1_combout ),
	.cout());
defparam \av_ld_byte2_data[7]~1 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[7]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte2_data[6]~2 (
	.dataa(src_data_22),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[6]~2_combout ),
	.cout());
defparam \av_ld_byte2_data[6]~2 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[6]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte2_data[5]~3 (
	.dataa(src_data_21),
	.datab(\av_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte2_data[5]~3_combout ),
	.cout());
defparam \av_ld_byte2_data[5]~3 .lut_mask = 16'hAACC;
defparam \av_ld_byte2_data[5]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[31]~16 (
	.dataa(\Add1~96_combout ),
	.datab(\E_logic_result[31]~14_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[31]~16_combout ),
	.cout());
defparam \W_alu_result[31]~16 .lut_mask = 16'hAACC;
defparam \W_alu_result[31]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[16]~17 (
	.dataa(\Add1~66_combout ),
	.datab(\E_logic_result[16]~17_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[16]~17_combout ),
	.cout());
defparam \W_alu_result[16]~17 .lut_mask = 16'hAACC;
defparam \W_alu_result[16]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[30]~18 (
	.dataa(\Add1~94_combout ),
	.datab(\E_logic_result[30]~18_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[30]~18_combout ),
	.cout());
defparam \W_alu_result[30]~18 .lut_mask = 16'hAACC;
defparam \W_alu_result[30]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[29]~19 (
	.dataa(\Add1~92_combout ),
	.datab(\E_logic_result[29]~19_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[29]~19_combout ),
	.cout());
defparam \W_alu_result[29]~19 .lut_mask = 16'hAACC;
defparam \W_alu_result[29]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[28]~20 (
	.dataa(\Add1~90_combout ),
	.datab(\E_logic_result[28]~20_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[28]~20_combout ),
	.cout());
defparam \W_alu_result[28]~20 .lut_mask = 16'hAACC;
defparam \W_alu_result[28]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[27]~21 (
	.dataa(\Add1~88_combout ),
	.datab(\E_logic_result[27]~21_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[27]~21_combout ),
	.cout());
defparam \W_alu_result[27]~21 .lut_mask = 16'hAACC;
defparam \W_alu_result[27]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[26]~22 (
	.dataa(\Add1~86_combout ),
	.datab(\E_logic_result[26]~22_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[26]~22_combout ),
	.cout());
defparam \W_alu_result[26]~22 .lut_mask = 16'hAACC;
defparam \W_alu_result[26]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[25]~23 (
	.dataa(\Add1~84_combout ),
	.datab(\E_logic_result[25]~23_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[25]~23_combout ),
	.cout());
defparam \W_alu_result[25]~23 .lut_mask = 16'hAACC;
defparam \W_alu_result[25]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[24]~24 (
	.dataa(\Add1~82_combout ),
	.datab(\E_logic_result[24]~24_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[24]~24_combout ),
	.cout());
defparam \W_alu_result[24]~24 .lut_mask = 16'hAACC;
defparam \W_alu_result[24]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[23]~25 (
	.dataa(\Add1~80_combout ),
	.datab(\E_logic_result[23]~25_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[23]~25_combout ),
	.cout());
defparam \W_alu_result[23]~25 .lut_mask = 16'hAACC;
defparam \W_alu_result[23]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[22]~26 (
	.dataa(\Add1~78_combout ),
	.datab(\E_logic_result[22]~26_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[22]~26_combout ),
	.cout());
defparam \W_alu_result[22]~26 .lut_mask = 16'hAACC;
defparam \W_alu_result[22]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[21]~27 (
	.dataa(\Add1~76_combout ),
	.datab(\E_logic_result[21]~27_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[21]~27_combout ),
	.cout());
defparam \W_alu_result[21]~27 .lut_mask = 16'hAACC;
defparam \W_alu_result[21]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[20]~28 (
	.dataa(\Add1~74_combout ),
	.datab(\E_logic_result[20]~28_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[20]~28_combout ),
	.cout());
defparam \W_alu_result[20]~28 .lut_mask = 16'hAACC;
defparam \W_alu_result[20]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[19]~29 (
	.dataa(\Add1~72_combout ),
	.datab(\E_logic_result[19]~29_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[19]~29_combout ),
	.cout());
defparam \W_alu_result[19]~29 .lut_mask = 16'hAACC;
defparam \W_alu_result[19]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[18]~30 (
	.dataa(\Add1~70_combout ),
	.datab(\E_logic_result[18]~30_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[18]~30_combout ),
	.cout());
defparam \W_alu_result[18]~30 .lut_mask = 16'hAACC;
defparam \W_alu_result[18]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[17]~31 (
	.dataa(\Add1~68_combout ),
	.datab(\E_logic_result[17]~31_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[17]~31_combout ),
	.cout());
defparam \W_alu_result[17]~31 .lut_mask = 16'hAACC;
defparam \W_alu_result[17]~31 .sum_lutc_input = "datac";

dffeas R_wr_dst_reg(
	.clk(clk_clk),
	.d(\D_wr_dst_reg~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_wr_dst_reg~q ),
	.prn(vcc));
defparam R_wr_dst_reg.is_wysiwyg = "true";
defparam R_wr_dst_reg.power_up = "low";

cycloneive_lcell_comb W_rf_wren(
	.dataa(r_sync_rst),
	.datab(\R_wr_dst_reg~q ),
	.datac(\W_valid~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\W_rf_wren~combout ),
	.cout());
defparam W_rf_wren.lut_mask = 16'hFEFE;
defparam W_rf_wren.sum_lutc_input = "datac";

dffeas \av_ld_byte0_data[0] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data_nxt[0]~40_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[7]~0_combout ),
	.q(\av_ld_byte0_data[0]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[0] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[0] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[0]~0 (
	.dataa(\R_ctrl_br_cmp~q ),
	.datab(\W_cmp_result~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\W_rf_wr_data[0]~0_combout ),
	.cout());
defparam \W_rf_wr_data[0]~0 .lut_mask = 16'hEEEE;
defparam \W_rf_wr_data[0]~0 .sum_lutc_input = "datac";

dffeas \W_control_rd_data[0] (
	.clk(clk_clk),
	.d(\E_control_rd_data[0]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_control_rd_data[0]~q ),
	.prn(vcc));
defparam \W_control_rd_data[0] .is_wysiwyg = "true";
defparam \W_control_rd_data[0] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[0]~1 (
	.dataa(\W_control_rd_data[0]~q ),
	.datab(\W_alu_result[0]~q ),
	.datac(\R_ctrl_rd_ctl_reg~q ),
	.datad(\R_ctrl_br_cmp~q ),
	.cin(gnd),
	.combout(\W_rf_wr_data[0]~1_combout ),
	.cout());
defparam \W_rf_wr_data[0]~1 .lut_mask = 16'hACFF;
defparam \W_rf_wr_data[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[0]~2 (
	.dataa(\av_ld_byte0_data[0]~q ),
	.datab(\W_rf_wr_data[0]~0_combout ),
	.datac(\W_rf_wr_data[0]~1_combout ),
	.datad(\R_ctrl_ld~q ),
	.cin(gnd),
	.combout(\W_rf_wr_data[0]~2_combout ),
	.cout());
defparam \W_rf_wr_data[0]~2 .lut_mask = 16'hFAFC;
defparam \W_rf_wr_data[0]~2 .sum_lutc_input = "datac";

dffeas \R_dst_regnum[0] (
	.clk(clk_clk),
	.d(\D_dst_regnum[0]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_dst_regnum[0]~q ),
	.prn(vcc));
defparam \R_dst_regnum[0] .is_wysiwyg = "true";
defparam \R_dst_regnum[0] .power_up = "low";

dffeas \R_dst_regnum[1] (
	.clk(clk_clk),
	.d(\D_dst_regnum[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_dst_regnum[1]~q ),
	.prn(vcc));
defparam \R_dst_regnum[1] .is_wysiwyg = "true";
defparam \R_dst_regnum[1] .power_up = "low";

dffeas \R_dst_regnum[2] (
	.clk(clk_clk),
	.d(\D_dst_regnum[2]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_dst_regnum[2]~q ),
	.prn(vcc));
defparam \R_dst_regnum[2] .is_wysiwyg = "true";
defparam \R_dst_regnum[2] .power_up = "low";

dffeas \R_dst_regnum[3] (
	.clk(clk_clk),
	.d(\D_dst_regnum[3]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_dst_regnum[3]~q ),
	.prn(vcc));
defparam \R_dst_regnum[3] .is_wysiwyg = "true";
defparam \R_dst_regnum[3] .power_up = "low";

dffeas \R_dst_regnum[4] (
	.clk(clk_clk),
	.d(\D_dst_regnum[4]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_dst_regnum[4]~q ),
	.prn(vcc));
defparam \R_dst_regnum[4] .is_wysiwyg = "true";
defparam \R_dst_regnum[4] .power_up = "low";

dffeas \D_iw[22] (
	.clk(clk_clk),
	.d(\F_iw[22]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[22]~q ),
	.prn(vcc));
defparam \D_iw[22] .is_wysiwyg = "true";
defparam \D_iw[22] .power_up = "low";

dffeas \D_iw[23] (
	.clk(clk_clk),
	.d(\F_iw[23]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[23]~q ),
	.prn(vcc));
defparam \D_iw[23] .is_wysiwyg = "true";
defparam \D_iw[23] .power_up = "low";

dffeas \D_iw[24] (
	.clk(clk_clk),
	.d(\F_iw[24]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[24]~q ),
	.prn(vcc));
defparam \D_iw[24] .is_wysiwyg = "true";
defparam \D_iw[24] .power_up = "low";

dffeas \D_iw[25] (
	.clk(clk_clk),
	.d(\F_iw[25]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[25]~q ),
	.prn(vcc));
defparam \D_iw[25] .is_wysiwyg = "true";
defparam \D_iw[25] .power_up = "low";

dffeas \D_iw[26] (
	.clk(clk_clk),
	.d(\F_iw[26]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[26]~q ),
	.prn(vcc));
defparam \D_iw[26] .is_wysiwyg = "true";
defparam \D_iw[26] .power_up = "low";

dffeas \av_ld_byte0_data[1] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data_nxt[1]~41_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[7]~0_combout ),
	.q(\av_ld_byte0_data[1]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[1] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[1] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[1]~3 (
	.dataa(\av_ld_byte0_data[1]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[1]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[1]~3_combout ),
	.cout());
defparam \W_rf_wr_data[1]~3 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[1]~3 .sum_lutc_input = "datac";

dffeas \av_ld_byte0_data[2] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data_nxt[2]~42_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[7]~0_combout ),
	.q(\av_ld_byte0_data[2]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[2] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[2] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[2]~4 (
	.dataa(\av_ld_byte0_data[2]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_2),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[2]~4_combout ),
	.cout());
defparam \W_rf_wr_data[2]~4 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[2]~4 .sum_lutc_input = "datac";

dffeas \av_ld_byte0_data[3] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data_nxt[3]~43_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[7]~0_combout ),
	.q(\av_ld_byte0_data[3]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[3] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[3] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[3]~5 (
	.dataa(\av_ld_byte0_data[3]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_3),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[3]~5_combout ),
	.cout());
defparam \W_rf_wr_data[3]~5 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[3]~5 .sum_lutc_input = "datac";

dffeas \av_ld_byte0_data[4] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data_nxt[4]~44_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[7]~0_combout ),
	.q(\av_ld_byte0_data[4]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[4] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[4] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[4]~6 (
	.dataa(\av_ld_byte0_data[4]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_4),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[4]~6_combout ),
	.cout());
defparam \W_rf_wr_data[4]~6 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[4]~6 .sum_lutc_input = "datac";

dffeas \av_ld_byte0_data[5] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data_nxt[5]~45_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[7]~0_combout ),
	.q(\av_ld_byte0_data[5]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[5] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[5] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[5]~7 (
	.dataa(\av_ld_byte0_data[5]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_5),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[5]~7_combout ),
	.cout());
defparam \W_rf_wr_data[5]~7 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[5]~7 .sum_lutc_input = "datac";

dffeas \av_ld_byte0_data[6] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data_nxt[6]~46_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[7]~0_combout ),
	.q(\av_ld_byte0_data[6]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[6] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[6] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[6]~8 (
	.dataa(\av_ld_byte0_data[6]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_6),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[6]~8_combout ),
	.cout());
defparam \W_rf_wr_data[6]~8 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[6]~8 .sum_lutc_input = "datac";

dffeas \av_ld_byte0_data[7] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data_nxt[7]~47_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\av_ld_byte0_data[7]~0_combout ),
	.q(\av_ld_byte0_data[7]~q ),
	.prn(vcc));
defparam \av_ld_byte0_data[7] .is_wysiwyg = "true";
defparam \av_ld_byte0_data[7] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[7]~9 (
	.dataa(\av_ld_byte0_data[7]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_7),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[7]~9_combout ),
	.cout());
defparam \W_rf_wr_data[7]~9 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[7]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_wr_dst_reg~0 (
	.dataa(\Equal0~11_combout ),
	.datab(\Equal0~12_combout ),
	.datac(\D_iw[5]~q ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_wr_dst_reg~0_combout ),
	.cout());
defparam \D_wr_dst_reg~0 .lut_mask = 16'hEFFF;
defparam \D_wr_dst_reg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_wr_dst_reg~1 (
	.dataa(\Equal0~13_combout ),
	.datab(\D_iw[1]~q ),
	.datac(\D_iw[2]~q ),
	.datad(\R_ctrl_br_nxt~0_combout ),
	.cin(gnd),
	.combout(\D_wr_dst_reg~1_combout ),
	.cout());
defparam \D_wr_dst_reg~1 .lut_mask = 16'hFEFF;
defparam \D_wr_dst_reg~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~14 (
	.dataa(\Equal0~4_combout ),
	.datab(gnd),
	.datac(\D_iw[5]~q ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\Equal0~14_combout ),
	.cout());
defparam \Equal0~14 .lut_mask = 16'hAFFF;
defparam \Equal0~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_implicit_dst_eretaddr~14 (
	.dataa(\Equal62~8_combout ),
	.datab(\Equal62~13_combout ),
	.datac(\D_iw[14]~q ),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~14_combout ),
	.cout());
defparam \D_ctrl_implicit_dst_eretaddr~14 .lut_mask = 16'hEFFE;
defparam \D_ctrl_implicit_dst_eretaddr~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_implicit_dst_eretaddr~15 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[12]~q ),
	.datac(\D_iw[13]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~15_combout ),
	.cout());
defparam \D_ctrl_implicit_dst_eretaddr~15 .lut_mask = 16'hFBFF;
defparam \D_ctrl_implicit_dst_eretaddr~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_implicit_dst_eretaddr~17 (
	.dataa(\Equal0~7_combout ),
	.datab(\D_ctrl_implicit_dst_eretaddr~14_combout ),
	.datac(\D_ctrl_implicit_dst_eretaddr~15_combout ),
	.datad(\D_ctrl_implicit_dst_eretaddr~16_combout ),
	.cin(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~17_combout ),
	.cout());
defparam \D_ctrl_implicit_dst_eretaddr~17 .lut_mask = 16'hFFFE;
defparam \D_ctrl_implicit_dst_eretaddr~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[1]~0 (
	.dataa(\D_iw[23]~q ),
	.datab(\D_iw[18]~q ),
	.datac(\D_ctrl_b_is_dst~2_combout ),
	.datad(\D_ctrl_implicit_dst_eretaddr~17_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[1]~0_combout ),
	.cout());
defparam \D_dst_regnum[1]~0 .lut_mask = 16'hACFF;
defparam \D_dst_regnum[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[1]~1 (
	.dataa(\Equal0~14_combout ),
	.datab(\D_ctrl_implicit_dst_eretaddr~13_combout ),
	.datac(\D_ctrl_exception~2_combout ),
	.datad(\D_dst_regnum[1]~0_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[1]~1_combout ),
	.cout());
defparam \D_dst_regnum[1]~1 .lut_mask = 16'hFFFE;
defparam \D_dst_regnum[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[4]~2 (
	.dataa(\D_iw[26]~q ),
	.datab(\D_iw[21]~q ),
	.datac(\D_ctrl_b_is_dst~2_combout ),
	.datad(\Equal0~14_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[4]~2_combout ),
	.cout());
defparam \D_dst_regnum[4]~2 .lut_mask = 16'hFFAC;
defparam \D_dst_regnum[4]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[4]~3 (
	.dataa(\D_ctrl_implicit_dst_eretaddr~13_combout ),
	.datab(\D_ctrl_exception~2_combout ),
	.datac(\D_ctrl_implicit_dst_eretaddr~17_combout ),
	.datad(\D_dst_regnum[4]~2_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[4]~3_combout ),
	.cout());
defparam \D_dst_regnum[4]~3 .lut_mask = 16'hFFF7;
defparam \D_dst_regnum[4]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[3]~4 (
	.dataa(\D_iw[25]~q ),
	.datab(\D_iw[20]~q ),
	.datac(\D_ctrl_b_is_dst~2_combout ),
	.datad(\Equal0~14_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[3]~4_combout ),
	.cout());
defparam \D_dst_regnum[3]~4 .lut_mask = 16'hFFAC;
defparam \D_dst_regnum[3]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[3]~5 (
	.dataa(\D_ctrl_implicit_dst_eretaddr~13_combout ),
	.datab(\D_ctrl_exception~2_combout ),
	.datac(\D_ctrl_implicit_dst_eretaddr~17_combout ),
	.datad(\D_dst_regnum[3]~4_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[3]~5_combout ),
	.cout());
defparam \D_dst_regnum[3]~5 .lut_mask = 16'hFFF7;
defparam \D_dst_regnum[3]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[4]~6 (
	.dataa(\Equal0~14_combout ),
	.datab(\D_ctrl_implicit_dst_eretaddr~17_combout ),
	.datac(\D_ctrl_implicit_dst_eretaddr~10_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_dst_regnum[4]~6_combout ),
	.cout());
defparam \D_dst_regnum[4]~6 .lut_mask = 16'hF7F7;
defparam \D_dst_regnum[4]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[4]~7 (
	.dataa(\D_ctrl_exception~2_combout ),
	.datab(\D_ctrl_implicit_dst_eretaddr~5_combout ),
	.datac(\D_ctrl_implicit_dst_eretaddr~12_combout ),
	.datad(\D_dst_regnum[4]~6_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[4]~7_combout ),
	.cout());
defparam \D_dst_regnum[4]~7 .lut_mask = 16'hFFFE;
defparam \D_dst_regnum[4]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[2]~8 (
	.dataa(\D_iw[24]~q ),
	.datab(\D_iw[19]~q ),
	.datac(\D_ctrl_b_is_dst~2_combout ),
	.datad(\D_dst_regnum[4]~7_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[2]~8_combout ),
	.cout());
defparam \D_dst_regnum[2]~8 .lut_mask = 16'hACFF;
defparam \D_dst_regnum[2]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~18 (
	.dataa(\D_dst_regnum[1]~1_combout ),
	.datab(\D_dst_regnum[4]~3_combout ),
	.datac(\D_dst_regnum[3]~5_combout ),
	.datad(\D_dst_regnum[2]~8_combout ),
	.cin(gnd),
	.combout(\Equal0~18_combout ),
	.cout());
defparam \Equal0~18 .lut_mask = 16'h7FFF;
defparam \Equal0~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_dst_regnum[0]~9 (
	.dataa(\D_iw[22]~q ),
	.datab(\D_iw[17]~q ),
	.datac(\D_ctrl_b_is_dst~2_combout ),
	.datad(\D_dst_regnum[4]~7_combout ),
	.cin(gnd),
	.combout(\D_dst_regnum[0]~9_combout ),
	.cout());
defparam \D_dst_regnum[0]~9 .lut_mask = 16'hACFF;
defparam \D_dst_regnum[0]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_wr_dst_reg~2 (
	.dataa(\D_wr_dst_reg~0_combout ),
	.datab(\D_wr_dst_reg~1_combout ),
	.datac(\Equal0~18_combout ),
	.datad(\D_dst_regnum[0]~9_combout ),
	.cin(gnd),
	.combout(\D_wr_dst_reg~2_combout ),
	.cout());
defparam \D_wr_dst_reg~2 .lut_mask = 16'hFF7F;
defparam \D_wr_dst_reg~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[0]~16 (
	.dataa(read_latency_shift_reg_02),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_0),
	.datad(av_readdata_pre_01),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[0]~16_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[0]~16 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[0]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[0]~17 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_04),
	.datac(q_b_0),
	.datad(av_readdata_pre_02),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[0]~17_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[0]~17 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[0]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[0]~18 (
	.dataa(\av_ld_byte0_data_nxt[0]~16_combout ),
	.datab(\av_ld_byte0_data_nxt[0]~17_combout ),
	.datac(src0_valid),
	.datad(av_readdata_pre_03),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[0]~18_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[0]~18 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[0]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_rshift8~0 (
	.dataa(\W_alu_result[1]~q ),
	.datab(\W_alu_result[0]~q ),
	.datac(\av_ld_align_cycle[0]~q ),
	.datad(\av_ld_align_cycle[1]~q ),
	.cin(gnd),
	.combout(\av_ld_rshift8~0_combout ),
	.cout());
defparam \av_ld_rshift8~0 .lut_mask = 16'hEFFF;
defparam \av_ld_rshift8~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_rshift8~1 (
	.dataa(\av_ld_aligning_data~q ),
	.datab(\av_ld_rshift8~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\av_ld_rshift8~1_combout ),
	.cout());
defparam \av_ld_rshift8~1 .lut_mask = 16'hEEEE;
defparam \av_ld_rshift8~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data[7]~0 (
	.dataa(\av_ld_aligning_data~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\av_ld_rshift8~0_combout ),
	.cin(gnd),
	.combout(\av_ld_byte0_data[7]~0_combout ),
	.cout());
defparam \av_ld_byte0_data[7]~0 .lut_mask = 16'hFF55;
defparam \av_ld_byte0_data[7]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_control_rd_data[0]~0 (
	.dataa(\D_iw[7]~q ),
	.datab(\W_ienable_reg[0]~q ),
	.datac(\W_bstatus_reg~q ),
	.datad(\D_iw[6]~q ),
	.cin(gnd),
	.combout(\E_control_rd_data[0]~0_combout ),
	.cout());
defparam \E_control_rd_data[0]~0 .lut_mask = 16'hFDFE;
defparam \E_control_rd_data[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_control_rd_data[0]~1 (
	.dataa(\D_iw[8]~q ),
	.datab(\W_ipending_reg[0]~q ),
	.datac(\D_iw[10]~q ),
	.datad(\D_iw[9]~q ),
	.cin(gnd),
	.combout(\E_control_rd_data[0]~1_combout ),
	.cout());
defparam \E_control_rd_data[0]~1 .lut_mask = 16'hEDDE;
defparam \E_control_rd_data[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_control_rd_data[0]~2 (
	.dataa(\W_status_reg_pie~q ),
	.datab(\D_iw[8]~q ),
	.datac(\E_control_rd_data[0]~1_combout ),
	.datad(\E_control_rd_data[0]~0_combout ),
	.cin(gnd),
	.combout(\E_control_rd_data[0]~2_combout ),
	.cout());
defparam \E_control_rd_data[0]~2 .lut_mask = 16'hEBBE;
defparam \E_control_rd_data[0]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_control_rd_data[0]~3 (
	.dataa(\W_estatus_reg~q ),
	.datab(\D_iw[7]~q ),
	.datac(\E_control_rd_data[0]~0_combout ),
	.datad(\E_control_rd_data[0]~2_combout ),
	.cin(gnd),
	.combout(\E_control_rd_data[0]~3_combout ),
	.cout());
defparam \E_control_rd_data[0]~3 .lut_mask = 16'hEBBE;
defparam \E_control_rd_data[0]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_ld_signed~1 (
	.dataa(\D_iw[2]~q ),
	.datab(\D_ctrl_ld_signed~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_ld_signed~1_combout ),
	.cout());
defparam \D_ctrl_ld_signed~1 .lut_mask = 16'hEEEE;
defparam \D_ctrl_ld_signed~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[22]~0 (
	.dataa(read_latency_shift_reg_01),
	.datab(mem_73_0),
	.datac(mem_55_0),
	.datad(av_readdata_pre_22),
	.cin(gnd),
	.combout(\F_iw[22]~0_combout ),
	.cout());
defparam \F_iw[22]~0 .lut_mask = 16'hFFFE;
defparam \F_iw[22]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[22]~1 (
	.dataa(\D_iw[27]~0_combout ),
	.datab(\F_iw[22]~0_combout ),
	.datac(q_a_22),
	.datad(read_latency_shift_reg_05),
	.cin(gnd),
	.combout(\F_iw[22]~1_combout ),
	.cout());
defparam \F_iw[22]~1 .lut_mask = 16'hFFFE;
defparam \F_iw[22]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[23]~2 (
	.dataa(read_latency_shift_reg_01),
	.datab(mem_73_0),
	.datac(mem_55_0),
	.datad(av_readdata_pre_23),
	.cin(gnd),
	.combout(\F_iw[23]~2_combout ),
	.cout());
defparam \F_iw[23]~2 .lut_mask = 16'hFFFE;
defparam \F_iw[23]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[23]~3 (
	.dataa(\D_iw[27]~0_combout ),
	.datab(\F_iw[23]~2_combout ),
	.datac(read_latency_shift_reg_05),
	.datad(q_a_23),
	.cin(gnd),
	.combout(\F_iw[23]~3_combout ),
	.cout());
defparam \F_iw[23]~3 .lut_mask = 16'hFFFE;
defparam \F_iw[23]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[24]~4 (
	.dataa(read_latency_shift_reg_01),
	.datab(mem_73_0),
	.datac(mem_55_0),
	.datad(av_readdata_pre_24),
	.cin(gnd),
	.combout(\F_iw[24]~4_combout ),
	.cout());
defparam \F_iw[24]~4 .lut_mask = 16'hFFFE;
defparam \F_iw[24]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[24]~5 (
	.dataa(\D_iw[27]~0_combout ),
	.datab(\F_iw[24]~4_combout ),
	.datac(read_latency_shift_reg_05),
	.datad(q_a_24),
	.cin(gnd),
	.combout(\F_iw[24]~5_combout ),
	.cout());
defparam \F_iw[24]~5 .lut_mask = 16'hFFFE;
defparam \F_iw[24]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[25]~6 (
	.dataa(read_latency_shift_reg_01),
	.datab(mem_73_0),
	.datac(mem_55_0),
	.datad(av_readdata_pre_25),
	.cin(gnd),
	.combout(\F_iw[25]~6_combout ),
	.cout());
defparam \F_iw[25]~6 .lut_mask = 16'hFFFE;
defparam \F_iw[25]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[25]~7 (
	.dataa(\D_iw[27]~0_combout ),
	.datab(\F_iw[25]~6_combout ),
	.datac(read_latency_shift_reg_05),
	.datad(q_a_25),
	.cin(gnd),
	.combout(\F_iw[25]~7_combout ),
	.cout());
defparam \F_iw[25]~7 .lut_mask = 16'hFFFE;
defparam \F_iw[25]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[26]~8 (
	.dataa(read_latency_shift_reg_01),
	.datab(mem_73_0),
	.datac(mem_55_0),
	.datad(av_readdata_pre_26),
	.cin(gnd),
	.combout(\F_iw[26]~8_combout ),
	.cout());
defparam \F_iw[26]~8 .lut_mask = 16'hFFFE;
defparam \F_iw[26]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[26]~9 (
	.dataa(\D_iw[27]~0_combout ),
	.datab(\F_iw[26]~8_combout ),
	.datac(read_latency_shift_reg_05),
	.datad(q_a_26),
	.cin(gnd),
	.combout(\F_iw[26]~9_combout ),
	.cout());
defparam \F_iw[26]~9 .lut_mask = 16'hFFFE;
defparam \F_iw[26]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[12]~10 (
	.dataa(\av_ld_byte1_data[4]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_12),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[12]~10_combout ),
	.cout());
defparam \W_rf_wr_data[12]~10 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[12]~10 .sum_lutc_input = "datac";

dffeas \D_iw[27] (
	.clk(clk_clk),
	.d(\F_iw[27]~44_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[27]~q ),
	.prn(vcc));
defparam \D_iw[27] .is_wysiwyg = "true";
defparam \D_iw[27] .power_up = "low";

dffeas \D_iw[28] (
	.clk(clk_clk),
	.d(\F_iw[28]~46_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[28]~q ),
	.prn(vcc));
defparam \D_iw[28] .is_wysiwyg = "true";
defparam \D_iw[28] .power_up = "low";

dffeas \D_iw[29] (
	.clk(clk_clk),
	.d(\F_iw[29]~48_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[29]~q ),
	.prn(vcc));
defparam \D_iw[29] .is_wysiwyg = "true";
defparam \D_iw[29] .power_up = "low";

dffeas \D_iw[30] (
	.clk(clk_clk),
	.d(\F_iw[30]~50_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[30]~q ),
	.prn(vcc));
defparam \D_iw[30] .is_wysiwyg = "true";
defparam \D_iw[30] .power_up = "low";

dffeas \D_iw[31] (
	.clk(clk_clk),
	.d(\F_iw[31]~52_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[31]~q ),
	.prn(vcc));
defparam \D_iw[31] .is_wysiwyg = "true";
defparam \D_iw[31] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[11]~11 (
	.dataa(\av_ld_byte1_data[3]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_11),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[11]~11_combout ),
	.cout());
defparam \W_rf_wr_data[11]~11 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[11]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[10]~12 (
	.dataa(\av_ld_byte1_data[2]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_10),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[10]~12_combout ),
	.cout());
defparam \W_rf_wr_data[10]~12 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[10]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[9]~13 (
	.dataa(\av_ld_byte1_data[1]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_9),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[9]~13_combout ),
	.cout());
defparam \W_rf_wr_data[9]~13 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[9]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[8]~14 (
	.dataa(\av_ld_byte1_data[0]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_8),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[8]~14_combout ),
	.cout());
defparam \W_rf_wr_data[8]~14 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[8]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[15]~15 (
	.dataa(\av_ld_byte1_data[7]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_15),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[15]~15_combout ),
	.cout());
defparam \W_rf_wr_data[15]~15 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[15]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[14]~16 (
	.dataa(\av_ld_byte1_data[6]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_14),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[14]~16_combout ),
	.cout());
defparam \W_rf_wr_data[14]~16 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[14]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[13]~17 (
	.dataa(\av_ld_byte1_data[5]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(W_alu_result_13),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[13]~17_combout ),
	.cout());
defparam \W_rf_wr_data[13]~17 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[13]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[1]~19 (
	.dataa(read_latency_shift_reg_02),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_110),
	.datad(av_readdata_pre_111),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[1]~19_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[1]~19 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[1]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[1]~20 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_04),
	.datac(q_b_1),
	.datad(av_readdata_pre_112),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[1]~20_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[1]~20 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[1]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[1]~21 (
	.dataa(\av_ld_byte0_data_nxt[1]~19_combout ),
	.datab(\av_ld_byte0_data_nxt[1]~20_combout ),
	.datac(src0_valid),
	.datad(av_readdata_pre_1),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[1]~21_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[1]~21 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[1]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[2]~22 (
	.dataa(read_latency_shift_reg_02),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_27),
	.datad(av_readdata_pre_28),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[2]~22_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[2]~22 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[2]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[2]~23 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_04),
	.datac(q_b_2),
	.datad(av_readdata_pre_29),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[2]~23_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[2]~23 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[2]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[2]~24 (
	.dataa(\av_ld_byte0_data_nxt[2]~22_combout ),
	.datab(\av_ld_byte0_data_nxt[2]~23_combout ),
	.datac(src0_valid),
	.datad(av_readdata_pre_2),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[2]~24_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[2]~24 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[2]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[3]~25 (
	.dataa(read_latency_shift_reg_02),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_31),
	.datad(av_readdata_pre_32),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[3]~25_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[3]~25 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[3]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[3]~26 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_04),
	.datac(q_b_3),
	.datad(av_readdata_pre_33),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[3]~26_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[3]~26 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[3]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[3]~27 (
	.dataa(\av_ld_byte0_data_nxt[3]~25_combout ),
	.datab(\av_ld_byte0_data_nxt[3]~26_combout ),
	.datac(src0_valid),
	.datad(av_readdata_pre_3),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[3]~27_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[3]~27 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[3]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[4]~28 (
	.dataa(read_latency_shift_reg_02),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_41),
	.datad(av_readdata_pre_42),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[4]~28_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[4]~28 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[4]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[4]~29 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_04),
	.datac(q_b_4),
	.datad(av_readdata_pre_43),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[4]~29_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[4]~29 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[4]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[4]~30 (
	.dataa(\av_ld_byte0_data_nxt[4]~28_combout ),
	.datab(\av_ld_byte0_data_nxt[4]~29_combout ),
	.datac(src0_valid),
	.datad(av_readdata_pre_4),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[4]~30_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[4]~30 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[4]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[5]~31 (
	.dataa(read_latency_shift_reg_02),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_51),
	.datad(av_readdata_pre_52),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[5]~31_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[5]~31 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[5]~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[5]~32 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_04),
	.datac(q_b_5),
	.datad(av_readdata_pre_53),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[5]~32_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[5]~32 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[5]~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[5]~33 (
	.dataa(\av_ld_byte0_data_nxt[5]~31_combout ),
	.datab(\av_ld_byte0_data_nxt[5]~32_combout ),
	.datac(src0_valid),
	.datad(av_readdata_pre_5),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[5]~33_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[5]~33 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[5]~33 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[6]~34 (
	.dataa(read_latency_shift_reg_02),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_61),
	.datad(av_readdata_pre_62),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[6]~34_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[6]~34 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[6]~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[6]~35 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_04),
	.datac(q_b_6),
	.datad(av_readdata_pre_63),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[6]~35_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[6]~35 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[6]~35 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[6]~36 (
	.dataa(\av_ld_byte0_data_nxt[6]~34_combout ),
	.datab(\av_ld_byte0_data_nxt[6]~35_combout ),
	.datac(src0_valid),
	.datad(av_readdata_pre_6),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[6]~36_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[6]~36 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[6]~36 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[7]~37 (
	.dataa(read_latency_shift_reg_02),
	.datab(read_latency_shift_reg_03),
	.datac(av_readdata_pre_71),
	.datad(av_readdata_pre_72),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[7]~37_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[7]~37 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[7]~37 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[7]~38 (
	.dataa(read_latency_shift_reg_0),
	.datab(read_latency_shift_reg_04),
	.datac(q_b_7),
	.datad(av_readdata_pre_73),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[7]~38_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[7]~38 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[7]~38 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[7]~39 (
	.dataa(\av_ld_byte0_data_nxt[7]~37_combout ),
	.datab(\av_ld_byte0_data_nxt[7]~38_combout ),
	.datac(src0_valid),
	.datad(av_readdata_pre_7),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[7]~39_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[7]~39 .lut_mask = 16'hFFFE;
defparam \av_ld_byte0_data_nxt[7]~39 .sum_lutc_input = "datac";

dffeas R_ctrl_ld_signed(
	.clk(clk_clk),
	.d(\D_ctrl_ld_signed~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_ld_signed~q ),
	.prn(vcc));
defparam R_ctrl_ld_signed.is_wysiwyg = "true";
defparam R_ctrl_ld_signed.power_up = "low";

cycloneive_lcell_comb \av_fill_bit~0 (
	.dataa(\R_ctrl_ld_signed~q ),
	.datab(\av_ld_byte1_data[7]~q ),
	.datac(\av_ld_byte0_data[7]~q ),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\av_fill_bit~0_combout ),
	.cout());
defparam \av_fill_bit~0 .lut_mask = 16'hFAFC;
defparam \av_fill_bit~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte1_data_en~0 (
	.dataa(\D_iw[4]~q ),
	.datab(\av_ld_rshift8~0_combout ),
	.datac(\av_ld_aligning_data~q ),
	.datad(\D_ctrl_mem16~0_combout ),
	.cin(gnd),
	.combout(\av_ld_byte1_data_en~0_combout ),
	.cout());
defparam \av_ld_byte1_data_en~0 .lut_mask = 16'hEFFF;
defparam \av_ld_byte1_data_en~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[27]~43 (
	.dataa(read_latency_shift_reg_01),
	.datab(mem_73_0),
	.datac(mem_55_0),
	.datad(av_readdata_pre_271),
	.cin(gnd),
	.combout(\F_iw[27]~43_combout ),
	.cout());
defparam \F_iw[27]~43 .lut_mask = 16'hFFFE;
defparam \F_iw[27]~43 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[27]~44 (
	.dataa(\D_iw[27]~0_combout ),
	.datab(\F_iw[27]~43_combout ),
	.datac(read_latency_shift_reg_05),
	.datad(q_a_27),
	.cin(gnd),
	.combout(\F_iw[27]~44_combout ),
	.cout());
defparam \F_iw[27]~44 .lut_mask = 16'hFFFE;
defparam \F_iw[27]~44 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[28]~45 (
	.dataa(read_latency_shift_reg_01),
	.datab(mem_73_0),
	.datac(mem_55_0),
	.datad(av_readdata_pre_281),
	.cin(gnd),
	.combout(\F_iw[28]~45_combout ),
	.cout());
defparam \F_iw[28]~45 .lut_mask = 16'hFFFE;
defparam \F_iw[28]~45 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[28]~46 (
	.dataa(\D_iw[27]~0_combout ),
	.datab(\F_iw[28]~45_combout ),
	.datac(read_latency_shift_reg_05),
	.datad(q_a_28),
	.cin(gnd),
	.combout(\F_iw[28]~46_combout ),
	.cout());
defparam \F_iw[28]~46 .lut_mask = 16'hFFFE;
defparam \F_iw[28]~46 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[29]~47 (
	.dataa(read_latency_shift_reg_01),
	.datab(mem_73_0),
	.datac(mem_55_0),
	.datad(av_readdata_pre_291),
	.cin(gnd),
	.combout(\F_iw[29]~47_combout ),
	.cout());
defparam \F_iw[29]~47 .lut_mask = 16'hFFFE;
defparam \F_iw[29]~47 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[29]~48 (
	.dataa(\D_iw[27]~0_combout ),
	.datab(\F_iw[29]~47_combout ),
	.datac(read_latency_shift_reg_05),
	.datad(q_a_29),
	.cin(gnd),
	.combout(\F_iw[29]~48_combout ),
	.cout());
defparam \F_iw[29]~48 .lut_mask = 16'hFFFE;
defparam \F_iw[29]~48 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[30]~49 (
	.dataa(read_latency_shift_reg_01),
	.datab(mem_73_0),
	.datac(mem_55_0),
	.datad(av_readdata_pre_30),
	.cin(gnd),
	.combout(\F_iw[30]~49_combout ),
	.cout());
defparam \F_iw[30]~49 .lut_mask = 16'hFFFE;
defparam \F_iw[30]~49 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[30]~50 (
	.dataa(\D_iw[27]~0_combout ),
	.datab(\F_iw[30]~49_combout ),
	.datac(read_latency_shift_reg_05),
	.datad(q_a_30),
	.cin(gnd),
	.combout(\F_iw[30]~50_combout ),
	.cout());
defparam \F_iw[30]~50 .lut_mask = 16'hFFFE;
defparam \F_iw[30]~50 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[31]~51 (
	.dataa(read_latency_shift_reg_01),
	.datab(mem_73_0),
	.datac(mem_55_0),
	.datad(av_readdata_pre_311),
	.cin(gnd),
	.combout(\F_iw[31]~51_combout ),
	.cout());
defparam \F_iw[31]~51 .lut_mask = 16'hFFFE;
defparam \F_iw[31]~51 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[31]~52 (
	.dataa(\D_iw[27]~0_combout ),
	.datab(\F_iw[31]~51_combout ),
	.datac(read_latency_shift_reg_05),
	.datad(q_a_31),
	.cin(gnd),
	.combout(\F_iw[31]~52_combout ),
	.cout());
defparam \F_iw[31]~52 .lut_mask = 16'hFFFE;
defparam \F_iw[31]~52 .sum_lutc_input = "datac";

dffeas \av_ld_byte3_data[0] (
	.clk(clk_clk),
	.d(\av_ld_byte3_data_nxt~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[0]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[0] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[0] .power_up = "low";

dffeas \av_ld_byte3_data[7] (
	.clk(clk_clk),
	.d(\av_ld_byte3_data_nxt~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[7]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[7] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[7] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[31]~18 (
	.dataa(\av_ld_byte3_data[7]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[31]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[31]~18_combout ),
	.cout());
defparam \W_rf_wr_data[31]~18 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[31]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[16]~19 (
	.dataa(\av_ld_byte2_data[0]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[16]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[16]~19_combout ),
	.cout());
defparam \W_rf_wr_data[16]~19 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[16]~19 .sum_lutc_input = "datac";

dffeas \av_ld_byte3_data[6] (
	.clk(clk_clk),
	.d(\av_ld_byte3_data_nxt~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[6]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[6] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[6] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[30]~20 (
	.dataa(\av_ld_byte3_data[6]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[30]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[30]~20_combout ),
	.cout());
defparam \W_rf_wr_data[30]~20 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[30]~20 .sum_lutc_input = "datac";

dffeas \av_ld_byte3_data[5] (
	.clk(clk_clk),
	.d(\av_ld_byte3_data_nxt~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[5]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[5] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[5] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[29]~21 (
	.dataa(\av_ld_byte3_data[5]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[29]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[29]~21_combout ),
	.cout());
defparam \W_rf_wr_data[29]~21 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[29]~21 .sum_lutc_input = "datac";

dffeas \av_ld_byte3_data[4] (
	.clk(clk_clk),
	.d(\av_ld_byte3_data_nxt~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[4]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[4] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[4] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[28]~22 (
	.dataa(\av_ld_byte3_data[4]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[28]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[28]~22_combout ),
	.cout());
defparam \W_rf_wr_data[28]~22 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[28]~22 .sum_lutc_input = "datac";

dffeas \av_ld_byte3_data[3] (
	.clk(clk_clk),
	.d(\av_ld_byte3_data_nxt~17_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[3]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[3] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[3] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[27]~23 (
	.dataa(\av_ld_byte3_data[3]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[27]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[27]~23_combout ),
	.cout());
defparam \W_rf_wr_data[27]~23 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[27]~23 .sum_lutc_input = "datac";

dffeas \av_ld_byte3_data[2] (
	.clk(clk_clk),
	.d(\av_ld_byte3_data_nxt~20_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[2]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[2] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[2] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[26]~24 (
	.dataa(\av_ld_byte3_data[2]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[26]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[26]~24_combout ),
	.cout());
defparam \W_rf_wr_data[26]~24 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[26]~24 .sum_lutc_input = "datac";

dffeas \av_ld_byte3_data[1] (
	.clk(clk_clk),
	.d(\av_ld_byte3_data_nxt~23_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\av_ld_rshift8~1_combout ),
	.q(\av_ld_byte3_data[1]~q ),
	.prn(vcc));
defparam \av_ld_byte3_data[1] .is_wysiwyg = "true";
defparam \av_ld_byte3_data[1] .power_up = "low";

cycloneive_lcell_comb \W_rf_wr_data[25]~25 (
	.dataa(\av_ld_byte3_data[1]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[25]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[25]~25_combout ),
	.cout());
defparam \W_rf_wr_data[25]~25 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[25]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[24]~26 (
	.dataa(\av_ld_byte3_data[0]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[24]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[24]~26_combout ),
	.cout());
defparam \W_rf_wr_data[24]~26 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[24]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[23]~27 (
	.dataa(\av_ld_byte2_data[7]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[23]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[23]~27_combout ),
	.cout());
defparam \W_rf_wr_data[23]~27 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[23]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[22]~28 (
	.dataa(\av_ld_byte2_data[6]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[22]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[22]~28_combout ),
	.cout());
defparam \W_rf_wr_data[22]~28 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[22]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[21]~29 (
	.dataa(\av_ld_byte2_data[5]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[21]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[21]~29_combout ),
	.cout());
defparam \W_rf_wr_data[21]~29 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[21]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[20]~30 (
	.dataa(\av_ld_byte2_data[4]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[20]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[20]~30_combout ),
	.cout());
defparam \W_rf_wr_data[20]~30 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[20]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[19]~31 (
	.dataa(\av_ld_byte2_data[3]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[19]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[19]~31_combout ),
	.cout());
defparam \W_rf_wr_data[19]~31 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[19]~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[18]~32 (
	.dataa(\av_ld_byte2_data[2]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[18]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[18]~32_combout ),
	.cout());
defparam \W_rf_wr_data[18]~32 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[18]~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_rf_wr_data[17]~33 (
	.dataa(\av_ld_byte2_data[1]~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\W_alu_result[17]~q ),
	.datad(\E_alu_result~0_combout ),
	.cin(gnd),
	.combout(\W_rf_wr_data[17]~33_combout ),
	.cout());
defparam \W_rf_wr_data[17]~33 .lut_mask = 16'hB8FF;
defparam \W_rf_wr_data[17]~33 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~0 (
	.dataa(read_latency_shift_reg_01),
	.datab(av_readdata_pre_24),
	.datac(mem_73_0),
	.datad(mem_55_0),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~0_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~0 .lut_mask = 16'hEFFF;
defparam \av_ld_byte3_data_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~1 (
	.dataa(read_latency_shift_reg_03),
	.datab(read_latency_shift_reg_04),
	.datac(q_b_24),
	.datad(av_readdata_pre_241),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~1_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~1 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~2 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(\av_ld_byte3_data_nxt~0_combout ),
	.datac(\av_ld_byte3_data_nxt~1_combout ),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~2_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~2 .lut_mask = 16'hFAFC;
defparam \av_ld_byte3_data_nxt~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~3 (
	.dataa(read_latency_shift_reg_01),
	.datab(av_readdata_pre_311),
	.datac(mem_73_0),
	.datad(mem_55_0),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~3_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~3 .lut_mask = 16'hEFFF;
defparam \av_ld_byte3_data_nxt~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~4 (
	.dataa(read_latency_shift_reg_03),
	.datab(read_latency_shift_reg_04),
	.datac(q_b_31),
	.datad(av_readdata_pre_312),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~4_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~4 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~5 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(\av_ld_byte3_data_nxt~3_combout ),
	.datac(\av_ld_byte3_data_nxt~4_combout ),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~5_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~5 .lut_mask = 16'hFAFC;
defparam \av_ld_byte3_data_nxt~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~6 (
	.dataa(read_latency_shift_reg_01),
	.datab(av_readdata_pre_30),
	.datac(mem_73_0),
	.datad(mem_55_0),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~6_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~6 .lut_mask = 16'hEFFF;
defparam \av_ld_byte3_data_nxt~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~7 (
	.dataa(read_latency_shift_reg_03),
	.datab(read_latency_shift_reg_04),
	.datac(q_b_30),
	.datad(av_readdata_pre_301),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~7_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~7 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~8 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(\av_ld_byte3_data_nxt~6_combout ),
	.datac(\av_ld_byte3_data_nxt~7_combout ),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~8_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~8 .lut_mask = 16'hFAFC;
defparam \av_ld_byte3_data_nxt~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~9 (
	.dataa(read_latency_shift_reg_01),
	.datab(av_readdata_pre_291),
	.datac(mem_73_0),
	.datad(mem_55_0),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~9_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~9 .lut_mask = 16'hEFFF;
defparam \av_ld_byte3_data_nxt~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~10 (
	.dataa(read_latency_shift_reg_03),
	.datab(read_latency_shift_reg_04),
	.datac(q_b_29),
	.datad(av_readdata_pre_292),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~10_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~10 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~11 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(\av_ld_byte3_data_nxt~9_combout ),
	.datac(\av_ld_byte3_data_nxt~10_combout ),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~11_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~11 .lut_mask = 16'hFAFC;
defparam \av_ld_byte3_data_nxt~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~12 (
	.dataa(read_latency_shift_reg_01),
	.datab(av_readdata_pre_281),
	.datac(mem_73_0),
	.datad(mem_55_0),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~12_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~12 .lut_mask = 16'hEFFF;
defparam \av_ld_byte3_data_nxt~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~13 (
	.dataa(read_latency_shift_reg_03),
	.datab(read_latency_shift_reg_04),
	.datac(q_b_28),
	.datad(av_readdata_pre_282),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~13_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~13 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~14 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(\av_ld_byte3_data_nxt~12_combout ),
	.datac(\av_ld_byte3_data_nxt~13_combout ),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~14_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~14 .lut_mask = 16'hFAFC;
defparam \av_ld_byte3_data_nxt~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~15 (
	.dataa(read_latency_shift_reg_01),
	.datab(av_readdata_pre_271),
	.datac(mem_73_0),
	.datad(mem_55_0),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~15_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~15 .lut_mask = 16'hEFFF;
defparam \av_ld_byte3_data_nxt~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~16 (
	.dataa(read_latency_shift_reg_03),
	.datab(read_latency_shift_reg_04),
	.datac(q_b_27),
	.datad(av_readdata_pre_272),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~16_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~16 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~17 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(\av_ld_byte3_data_nxt~15_combout ),
	.datac(\av_ld_byte3_data_nxt~16_combout ),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~17_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~17 .lut_mask = 16'hFAFC;
defparam \av_ld_byte3_data_nxt~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~18 (
	.dataa(read_latency_shift_reg_01),
	.datab(av_readdata_pre_26),
	.datac(mem_73_0),
	.datad(mem_55_0),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~18_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~18 .lut_mask = 16'hEFFF;
defparam \av_ld_byte3_data_nxt~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~19 (
	.dataa(read_latency_shift_reg_03),
	.datab(read_latency_shift_reg_04),
	.datac(q_b_26),
	.datad(av_readdata_pre_261),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~19_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~19 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~20 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(\av_ld_byte3_data_nxt~18_combout ),
	.datac(\av_ld_byte3_data_nxt~19_combout ),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~20_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~20 .lut_mask = 16'hFAFC;
defparam \av_ld_byte3_data_nxt~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~21 (
	.dataa(read_latency_shift_reg_01),
	.datab(av_readdata_pre_25),
	.datac(mem_73_0),
	.datad(mem_55_0),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~21_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~21 .lut_mask = 16'hEFFF;
defparam \av_ld_byte3_data_nxt~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~22 (
	.dataa(read_latency_shift_reg_03),
	.datab(read_latency_shift_reg_04),
	.datac(q_b_25),
	.datad(av_readdata_pre_251),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~22_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~22 .lut_mask = 16'hFFFE;
defparam \av_ld_byte3_data_nxt~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte3_data_nxt~23 (
	.dataa(\av_fill_bit~0_combout ),
	.datab(\av_ld_byte3_data_nxt~21_combout ),
	.datac(\av_ld_byte3_data_nxt~22_combout ),
	.datad(\av_ld_aligning_data~q ),
	.cin(gnd),
	.combout(\av_ld_byte3_data_nxt~23_combout ),
	.cout());
defparam \av_ld_byte3_data_nxt~23 .lut_mask = 16'hFAFC;
defparam \av_ld_byte3_data_nxt~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[0]~40 (
	.dataa(\av_ld_aligning_data~q ),
	.datab(\av_ld_rshift8~0_combout ),
	.datac(\av_ld_byte1_data[0]~q ),
	.datad(\av_ld_byte0_data_nxt[0]~18_combout ),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[0]~40_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[0]~40 .lut_mask = 16'hFFF6;
defparam \av_ld_byte0_data_nxt[0]~40 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[1]~41 (
	.dataa(\av_ld_aligning_data~q ),
	.datab(\av_ld_rshift8~0_combout ),
	.datac(\av_ld_byte1_data[1]~q ),
	.datad(\av_ld_byte0_data_nxt[1]~21_combout ),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[1]~41_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[1]~41 .lut_mask = 16'hFFF6;
defparam \av_ld_byte0_data_nxt[1]~41 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[2]~42 (
	.dataa(\av_ld_aligning_data~q ),
	.datab(\av_ld_rshift8~0_combout ),
	.datac(\av_ld_byte1_data[2]~q ),
	.datad(\av_ld_byte0_data_nxt[2]~24_combout ),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[2]~42_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[2]~42 .lut_mask = 16'hFFF6;
defparam \av_ld_byte0_data_nxt[2]~42 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[3]~43 (
	.dataa(\av_ld_aligning_data~q ),
	.datab(\av_ld_rshift8~0_combout ),
	.datac(\av_ld_byte1_data[3]~q ),
	.datad(\av_ld_byte0_data_nxt[3]~27_combout ),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[3]~43_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[3]~43 .lut_mask = 16'hFFF6;
defparam \av_ld_byte0_data_nxt[3]~43 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[4]~44 (
	.dataa(\av_ld_aligning_data~q ),
	.datab(\av_ld_rshift8~0_combout ),
	.datac(\av_ld_byte1_data[4]~q ),
	.datad(\av_ld_byte0_data_nxt[4]~30_combout ),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[4]~44_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[4]~44 .lut_mask = 16'hFFF6;
defparam \av_ld_byte0_data_nxt[4]~44 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[5]~45 (
	.dataa(\av_ld_aligning_data~q ),
	.datab(\av_ld_rshift8~0_combout ),
	.datac(\av_ld_byte1_data[5]~q ),
	.datad(\av_ld_byte0_data_nxt[5]~33_combout ),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[5]~45_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[5]~45 .lut_mask = 16'hFFF6;
defparam \av_ld_byte0_data_nxt[5]~45 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[6]~46 (
	.dataa(\av_ld_aligning_data~q ),
	.datab(\av_ld_rshift8~0_combout ),
	.datac(\av_ld_byte1_data[6]~q ),
	.datad(\av_ld_byte0_data_nxt[6]~36_combout ),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[6]~46_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[6]~46 .lut_mask = 16'hFFF6;
defparam \av_ld_byte0_data_nxt[6]~46 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_byte0_data_nxt[7]~47 (
	.dataa(\av_ld_aligning_data~q ),
	.datab(\av_ld_rshift8~0_combout ),
	.datac(\av_ld_byte1_data[7]~q ),
	.datad(\av_ld_byte0_data_nxt[7]~39_combout ),
	.cin(gnd),
	.combout(\av_ld_byte0_data_nxt[7]~47_combout ),
	.cout());
defparam \av_ld_byte0_data_nxt[7]~47 .lut_mask = 16'hFFF6;
defparam \av_ld_byte0_data_nxt[7]~47 .sum_lutc_input = "datac";

dffeas \W_alu_result[12] (
	.clk(clk_clk),
	.d(\W_alu_result[12]~3_combout ),
	.asdata(\E_shift_rot_result[12]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_12),
	.prn(vcc));
defparam \W_alu_result[12] .is_wysiwyg = "true";
defparam \W_alu_result[12] .power_up = "low";

dffeas \W_alu_result[15] (
	.clk(clk_clk),
	.d(\W_alu_result[15]~0_combout ),
	.asdata(\E_shift_rot_result[15]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_15),
	.prn(vcc));
defparam \W_alu_result[15] .is_wysiwyg = "true";
defparam \W_alu_result[15] .power_up = "low";

dffeas \W_alu_result[14] (
	.clk(clk_clk),
	.d(\W_alu_result[14]~1_combout ),
	.asdata(\E_shift_rot_result[14]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_14),
	.prn(vcc));
defparam \W_alu_result[14] .is_wysiwyg = "true";
defparam \W_alu_result[14] .power_up = "low";

dffeas \W_alu_result[13] (
	.clk(clk_clk),
	.d(\W_alu_result[13]~2_combout ),
	.asdata(\E_shift_rot_result[13]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_13),
	.prn(vcc));
defparam \W_alu_result[13] .is_wysiwyg = "true";
defparam \W_alu_result[13] .power_up = "low";

dffeas \W_alu_result[11] (
	.clk(clk_clk),
	.d(\W_alu_result[11]~4_combout ),
	.asdata(\E_shift_rot_result[11]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_11),
	.prn(vcc));
defparam \W_alu_result[11] .is_wysiwyg = "true";
defparam \W_alu_result[11] .power_up = "low";

dffeas \W_alu_result[10] (
	.clk(clk_clk),
	.d(\W_alu_result[10]~5_combout ),
	.asdata(\E_shift_rot_result[10]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_10),
	.prn(vcc));
defparam \W_alu_result[10] .is_wysiwyg = "true";
defparam \W_alu_result[10] .power_up = "low";

dffeas \W_alu_result[9] (
	.clk(clk_clk),
	.d(\W_alu_result[9]~6_combout ),
	.asdata(\E_shift_rot_result[9]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_9),
	.prn(vcc));
defparam \W_alu_result[9] .is_wysiwyg = "true";
defparam \W_alu_result[9] .power_up = "low";

dffeas \W_alu_result[8] (
	.clk(clk_clk),
	.d(\W_alu_result[8]~7_combout ),
	.asdata(\E_shift_rot_result[8]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_8),
	.prn(vcc));
defparam \W_alu_result[8] .is_wysiwyg = "true";
defparam \W_alu_result[8] .power_up = "low";

dffeas \W_alu_result[7] (
	.clk(clk_clk),
	.d(\W_alu_result[7]~8_combout ),
	.asdata(\E_shift_rot_result[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_7),
	.prn(vcc));
defparam \W_alu_result[7] .is_wysiwyg = "true";
defparam \W_alu_result[7] .power_up = "low";

dffeas \W_alu_result[6] (
	.clk(clk_clk),
	.d(\W_alu_result[6]~9_combout ),
	.asdata(\E_shift_rot_result[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_6),
	.prn(vcc));
defparam \W_alu_result[6] .is_wysiwyg = "true";
defparam \W_alu_result[6] .power_up = "low";

dffeas \W_alu_result[5] (
	.clk(clk_clk),
	.d(\W_alu_result[5]~10_combout ),
	.asdata(\E_shift_rot_result[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_5),
	.prn(vcc));
defparam \W_alu_result[5] .is_wysiwyg = "true";
defparam \W_alu_result[5] .power_up = "low";

dffeas \W_alu_result[4] (
	.clk(clk_clk),
	.d(\W_alu_result[4]~11_combout ),
	.asdata(\E_shift_rot_result[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_4),
	.prn(vcc));
defparam \W_alu_result[4] .is_wysiwyg = "true";
defparam \W_alu_result[4] .power_up = "low";

dffeas \W_alu_result[3] (
	.clk(clk_clk),
	.d(\W_alu_result[3]~12_combout ),
	.asdata(\E_shift_rot_result[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_3),
	.prn(vcc));
defparam \W_alu_result[3] .is_wysiwyg = "true";
defparam \W_alu_result[3] .power_up = "low";

dffeas \W_alu_result[2] (
	.clk(clk_clk),
	.d(\W_alu_result[2]~13_combout ),
	.asdata(\E_shift_rot_result[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\E_alu_result~0_combout ),
	.sload(\R_ctrl_shift_rot~q ),
	.ena(vcc),
	.q(W_alu_result_2),
	.prn(vcc));
defparam \W_alu_result[2] .is_wysiwyg = "true";
defparam \W_alu_result[2] .power_up = "low";

dffeas \d_writedata[24] (
	.clk(clk_clk),
	.d(\d_writedata[24]~0_combout ),
	.asdata(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_24),
	.prn(vcc));
defparam \d_writedata[24] .is_wysiwyg = "true";
defparam \d_writedata[24] .power_up = "low";

dffeas \d_writedata[25] (
	.clk(clk_clk),
	.d(\d_writedata[25]~1_combout ),
	.asdata(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_25),
	.prn(vcc));
defparam \d_writedata[25] .is_wysiwyg = "true";
defparam \d_writedata[25] .power_up = "low";

dffeas \d_writedata[26] (
	.clk(clk_clk),
	.d(\d_writedata[26]~2_combout ),
	.asdata(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_26),
	.prn(vcc));
defparam \d_writedata[26] .is_wysiwyg = "true";
defparam \d_writedata[26] .power_up = "low";

dffeas \d_writedata[27] (
	.clk(clk_clk),
	.d(\d_writedata[27]~3_combout ),
	.asdata(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_27),
	.prn(vcc));
defparam \d_writedata[27] .is_wysiwyg = "true";
defparam \d_writedata[27] .power_up = "low";

dffeas \d_writedata[28] (
	.clk(clk_clk),
	.d(\d_writedata[28]~4_combout ),
	.asdata(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_28),
	.prn(vcc));
defparam \d_writedata[28] .is_wysiwyg = "true";
defparam \d_writedata[28] .power_up = "low";

dffeas \d_writedata[29] (
	.clk(clk_clk),
	.d(\d_writedata[29]~5_combout ),
	.asdata(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_29),
	.prn(vcc));
defparam \d_writedata[29] .is_wysiwyg = "true";
defparam \d_writedata[29] .power_up = "low";

dffeas \d_writedata[30] (
	.clk(clk_clk),
	.d(\d_writedata[30]~6_combout ),
	.asdata(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_30),
	.prn(vcc));
defparam \d_writedata[30] .is_wysiwyg = "true";
defparam \d_writedata[30] .power_up = "low";

dffeas \d_writedata[31] (
	.clk(clk_clk),
	.d(\d_writedata[31]~7_combout ),
	.asdata(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_ctrl_mem8~1_combout ),
	.ena(vcc),
	.q(d_writedata_31),
	.prn(vcc));
defparam \d_writedata[31] .is_wysiwyg = "true";
defparam \d_writedata[31] .power_up = "low";

dffeas \d_writedata[0] (
	.clk(clk_clk),
	.d(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_0),
	.prn(vcc));
defparam \d_writedata[0] .is_wysiwyg = "true";
defparam \d_writedata[0] .power_up = "low";

dffeas d_write(
	.clk(clk_clk),
	.d(\E_st_stall~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_write1),
	.prn(vcc));
defparam d_write.is_wysiwyg = "true";
defparam d_write.power_up = "low";

dffeas \d_writedata[1] (
	.clk(clk_clk),
	.d(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_1),
	.prn(vcc));
defparam \d_writedata[1] .is_wysiwyg = "true";
defparam \d_writedata[1] .power_up = "low";

dffeas \d_writedata[2] (
	.clk(clk_clk),
	.d(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_2),
	.prn(vcc));
defparam \d_writedata[2] .is_wysiwyg = "true";
defparam \d_writedata[2] .power_up = "low";

dffeas \d_writedata[3] (
	.clk(clk_clk),
	.d(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_3),
	.prn(vcc));
defparam \d_writedata[3] .is_wysiwyg = "true";
defparam \d_writedata[3] .power_up = "low";

dffeas \d_writedata[4] (
	.clk(clk_clk),
	.d(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_4),
	.prn(vcc));
defparam \d_writedata[4] .is_wysiwyg = "true";
defparam \d_writedata[4] .power_up = "low";

dffeas \d_writedata[5] (
	.clk(clk_clk),
	.d(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_5),
	.prn(vcc));
defparam \d_writedata[5] .is_wysiwyg = "true";
defparam \d_writedata[5] .power_up = "low";

dffeas \d_writedata[6] (
	.clk(clk_clk),
	.d(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_6),
	.prn(vcc));
defparam \d_writedata[6] .is_wysiwyg = "true";
defparam \d_writedata[6] .power_up = "low";

dffeas \d_writedata[7] (
	.clk(clk_clk),
	.d(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_7),
	.prn(vcc));
defparam \d_writedata[7] .is_wysiwyg = "true";
defparam \d_writedata[7] .power_up = "low";

dffeas d_read(
	.clk(clk_clk),
	.d(\d_read_nxt~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_read1),
	.prn(vcc));
defparam d_read.is_wysiwyg = "true";
defparam d_read.power_up = "low";

dffeas \F_pc[10] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[10]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_10),
	.prn(vcc));
defparam \F_pc[10] .is_wysiwyg = "true";
defparam \F_pc[10] .power_up = "low";

dffeas \F_pc[9] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[9]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_9),
	.prn(vcc));
defparam \F_pc[9] .is_wysiwyg = "true";
defparam \F_pc[9] .power_up = "low";

dffeas \F_pc[8] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[8]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_8),
	.prn(vcc));
defparam \F_pc[8] .is_wysiwyg = "true";
defparam \F_pc[8] .power_up = "low";

dffeas \F_pc[7] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[7]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_7),
	.prn(vcc));
defparam \F_pc[7] .is_wysiwyg = "true";
defparam \F_pc[7] .power_up = "low";

dffeas \F_pc[6] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[6]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_6),
	.prn(vcc));
defparam \F_pc[6] .is_wysiwyg = "true";
defparam \F_pc[6] .power_up = "low";

dffeas \F_pc[5] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[5]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_5),
	.prn(vcc));
defparam \F_pc[5] .is_wysiwyg = "true";
defparam \F_pc[5] .power_up = "low";

dffeas \F_pc[4] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[4]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_4),
	.prn(vcc));
defparam \F_pc[4] .is_wysiwyg = "true";
defparam \F_pc[4] .power_up = "low";

dffeas \F_pc[3] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[3]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_3),
	.prn(vcc));
defparam \F_pc[3] .is_wysiwyg = "true";
defparam \F_pc[3] .power_up = "low";

dffeas \F_pc[2] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[2]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_2),
	.prn(vcc));
defparam \F_pc[2] .is_wysiwyg = "true";
defparam \F_pc[2] .power_up = "low";

dffeas \F_pc[1] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[1]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_1),
	.prn(vcc));
defparam \F_pc[1] .is_wysiwyg = "true";
defparam \F_pc[1] .power_up = "low";

dffeas \F_pc[0] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[0]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_0),
	.prn(vcc));
defparam \F_pc[0] .is_wysiwyg = "true";
defparam \F_pc[0] .power_up = "low";

dffeas \F_pc[13] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[13]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_13),
	.prn(vcc));
defparam \F_pc[13] .is_wysiwyg = "true";
defparam \F_pc[13] .power_up = "low";

dffeas \F_pc[12] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[12]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_12),
	.prn(vcc));
defparam \F_pc[12] .is_wysiwyg = "true";
defparam \F_pc[12] .power_up = "low";

dffeas \F_pc[11] (
	.clk(clk_clk),
	.d(\F_pc_no_crst_nxt[11]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_valid~q ),
	.q(F_pc_11),
	.prn(vcc));
defparam \F_pc[11] .is_wysiwyg = "true";
defparam \F_pc[11] .power_up = "low";

dffeas i_read(
	.clk(clk_clk),
	.d(\i_read_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(i_read1),
	.prn(vcc));
defparam i_read.is_wysiwyg = "true";
defparam i_read.power_up = "low";

dffeas hbreak_enabled(
	.clk(clk_clk),
	.d(\hbreak_enabled~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\E_valid_from_R~q ),
	.q(hbreak_enabled1),
	.prn(vcc));
defparam hbreak_enabled.is_wysiwyg = "true";
defparam hbreak_enabled.power_up = "low";

dffeas \d_byteenable[0] (
	.clk(clk_clk),
	.d(\E_mem_byte_en[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_byteenable_0),
	.prn(vcc));
defparam \d_byteenable[0] .is_wysiwyg = "true";
defparam \d_byteenable[0] .power_up = "low";

dffeas \d_writedata[22] (
	.clk(clk_clk),
	.d(\E_st_data[22]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_22),
	.prn(vcc));
defparam \d_writedata[22] .is_wysiwyg = "true";
defparam \d_writedata[22] .power_up = "low";

dffeas \d_byteenable[2] (
	.clk(clk_clk),
	.d(\E_mem_byte_en[2]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_byteenable_2),
	.prn(vcc));
defparam \d_byteenable[2] .is_wysiwyg = "true";
defparam \d_byteenable[2] .power_up = "low";

dffeas \d_writedata[23] (
	.clk(clk_clk),
	.d(\E_st_data[23]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_23),
	.prn(vcc));
defparam \d_writedata[23] .is_wysiwyg = "true";
defparam \d_writedata[23] .power_up = "low";

dffeas \d_byteenable[3] (
	.clk(clk_clk),
	.d(\E_mem_byte_en[3]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_byteenable_3),
	.prn(vcc));
defparam \d_byteenable[3] .is_wysiwyg = "true";
defparam \d_byteenable[3] .power_up = "low";

dffeas \d_writedata[11] (
	.clk(clk_clk),
	.d(\E_st_data[11]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_11),
	.prn(vcc));
defparam \d_writedata[11] .is_wysiwyg = "true";
defparam \d_writedata[11] .power_up = "low";

dffeas \d_byteenable[1] (
	.clk(clk_clk),
	.d(\E_mem_byte_en[1]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_byteenable_1),
	.prn(vcc));
defparam \d_byteenable[1] .is_wysiwyg = "true";
defparam \d_byteenable[1] .power_up = "low";

dffeas \d_writedata[13] (
	.clk(clk_clk),
	.d(\E_st_data[13]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_13),
	.prn(vcc));
defparam \d_writedata[13] .is_wysiwyg = "true";
defparam \d_writedata[13] .power_up = "low";

dffeas \d_writedata[16] (
	.clk(clk_clk),
	.d(\E_st_data[16]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_16),
	.prn(vcc));
defparam \d_writedata[16] .is_wysiwyg = "true";
defparam \d_writedata[16] .power_up = "low";

dffeas \d_writedata[12] (
	.clk(clk_clk),
	.d(\E_st_data[12]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_12),
	.prn(vcc));
defparam \d_writedata[12] .is_wysiwyg = "true";
defparam \d_writedata[12] .power_up = "low";

dffeas \d_writedata[14] (
	.clk(clk_clk),
	.d(\E_st_data[14]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_14),
	.prn(vcc));
defparam \d_writedata[14] .is_wysiwyg = "true";
defparam \d_writedata[14] .power_up = "low";

dffeas \d_writedata[15] (
	.clk(clk_clk),
	.d(\E_st_data[15]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_15),
	.prn(vcc));
defparam \d_writedata[15] .is_wysiwyg = "true";
defparam \d_writedata[15] .power_up = "low";

dffeas \d_writedata[18] (
	.clk(clk_clk),
	.d(\E_st_data[18]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_18),
	.prn(vcc));
defparam \d_writedata[18] .is_wysiwyg = "true";
defparam \d_writedata[18] .power_up = "low";

dffeas \d_writedata[17] (
	.clk(clk_clk),
	.d(\E_st_data[17]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_17),
	.prn(vcc));
defparam \d_writedata[17] .is_wysiwyg = "true";
defparam \d_writedata[17] .power_up = "low";

dffeas \d_writedata[10] (
	.clk(clk_clk),
	.d(\E_st_data[10]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_10),
	.prn(vcc));
defparam \d_writedata[10] .is_wysiwyg = "true";
defparam \d_writedata[10] .power_up = "low";

dffeas \d_writedata[9] (
	.clk(clk_clk),
	.d(\E_st_data[9]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_9),
	.prn(vcc));
defparam \d_writedata[9] .is_wysiwyg = "true";
defparam \d_writedata[9] .power_up = "low";

dffeas \d_writedata[8] (
	.clk(clk_clk),
	.d(\E_st_data[8]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_8),
	.prn(vcc));
defparam \d_writedata[8] .is_wysiwyg = "true";
defparam \d_writedata[8] .power_up = "low";

dffeas \d_writedata[21] (
	.clk(clk_clk),
	.d(\E_st_data[21]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_21),
	.prn(vcc));
defparam \d_writedata[21] .is_wysiwyg = "true";
defparam \d_writedata[21] .power_up = "low";

dffeas \d_writedata[19] (
	.clk(clk_clk),
	.d(\E_st_data[19]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_19),
	.prn(vcc));
defparam \d_writedata[19] .is_wysiwyg = "true";
defparam \d_writedata[19] .power_up = "low";

dffeas \d_writedata[20] (
	.clk(clk_clk),
	.d(\E_st_data[20]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_writedata_20),
	.prn(vcc));
defparam \d_writedata[20] .is_wysiwyg = "true";
defparam \d_writedata[20] .power_up = "low";

cycloneive_lcell_comb \F_valid~0 (
	.dataa(src1_valid),
	.datab(read_latency_shift_reg_05),
	.datac(gnd),
	.datad(i_read1),
	.cin(gnd),
	.combout(\F_valid~0_combout ),
	.cout());
defparam \F_valid~0 .lut_mask = 16'hEEFF;
defparam \F_valid~0 .sum_lutc_input = "datac";

dffeas D_valid(
	.clk(clk_clk),
	.d(\F_valid~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\D_valid~q ),
	.prn(vcc));
defparam D_valid.is_wysiwyg = "true";
defparam D_valid.power_up = "low";

dffeas R_valid(
	.clk(clk_clk),
	.d(\D_valid~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_valid~q ),
	.prn(vcc));
defparam R_valid.is_wysiwyg = "true";
defparam R_valid.power_up = "low";

cycloneive_lcell_comb \F_iw[1]~15 (
	.dataa(src_payload3),
	.datab(src1_valid),
	.datac(av_readdata_pre_1),
	.datad(\D_iw[27]~0_combout ),
	.cin(gnd),
	.combout(\F_iw[1]~15_combout ),
	.cout());
defparam \F_iw[1]~15 .lut_mask = 16'hFEFF;
defparam \F_iw[1]~15 .sum_lutc_input = "datac";

dffeas \D_iw[1] (
	.clk(clk_clk),
	.d(\F_iw[1]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[1]~q ),
	.prn(vcc));
defparam \D_iw[1] .is_wysiwyg = "true";
defparam \D_iw[1] .power_up = "low";

cycloneive_lcell_comb \F_iw[0]~16 (
	.dataa(read_latency_shift_reg_01),
	.datab(mem_73_0),
	.datac(mem_55_0),
	.datad(av_readdata_pre_03),
	.cin(gnd),
	.combout(\F_iw[0]~16_combout ),
	.cout());
defparam \F_iw[0]~16 .lut_mask = 16'hFFFE;
defparam \F_iw[0]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[0]~17 (
	.dataa(\D_iw[27]~0_combout ),
	.datab(\F_iw[0]~16_combout ),
	.datac(q_a_0),
	.datad(read_latency_shift_reg_05),
	.cin(gnd),
	.combout(\F_iw[0]~17_combout ),
	.cout());
defparam \F_iw[0]~17 .lut_mask = 16'hFFFE;
defparam \F_iw[0]~17 .sum_lutc_input = "datac";

dffeas \D_iw[0] (
	.clk(clk_clk),
	.d(\F_iw[0]~17_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[0]~q ),
	.prn(vcc));
defparam \D_iw[0] .is_wysiwyg = "true";
defparam \D_iw[0] .power_up = "low";

cycloneive_lcell_comb \F_iw[3]~18 (
	.dataa(src_payload4),
	.datab(src1_valid),
	.datac(av_readdata_pre_3),
	.datad(\D_iw[27]~0_combout ),
	.cin(gnd),
	.combout(\F_iw[3]~18_combout ),
	.cout());
defparam \F_iw[3]~18 .lut_mask = 16'hFEFF;
defparam \F_iw[3]~18 .sum_lutc_input = "datac";

dffeas \D_iw[3] (
	.clk(clk_clk),
	.d(\F_iw[3]~18_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[3]~q ),
	.prn(vcc));
defparam \D_iw[3] .is_wysiwyg = "true";
defparam \D_iw[3] .power_up = "low";

cycloneive_lcell_comb \F_iw[2]~19 (
	.dataa(read_latency_shift_reg_01),
	.datab(mem_73_0),
	.datac(mem_55_0),
	.datad(av_readdata_pre_2),
	.cin(gnd),
	.combout(\F_iw[2]~19_combout ),
	.cout());
defparam \F_iw[2]~19 .lut_mask = 16'hFFFE;
defparam \F_iw[2]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[2]~20 (
	.dataa(\D_iw[27]~0_combout ),
	.datab(\F_iw[2]~19_combout ),
	.datac(read_latency_shift_reg_05),
	.datad(q_a_2),
	.cin(gnd),
	.combout(\F_iw[2]~20_combout ),
	.cout());
defparam \F_iw[2]~20 .lut_mask = 16'hFFFE;
defparam \F_iw[2]~20 .sum_lutc_input = "datac";

dffeas \D_iw[2] (
	.clk(clk_clk),
	.d(\F_iw[2]~20_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[2]~q ),
	.prn(vcc));
defparam \D_iw[2] .is_wysiwyg = "true";
defparam \D_iw[2] .power_up = "low";

cycloneive_lcell_comb \Equal0~2 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~2_combout ),
	.cout());
defparam \Equal0~2 .lut_mask = 16'hFBFF;
defparam \Equal0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[5]~21 (
	.dataa(src_payload5),
	.datab(src1_valid),
	.datac(av_readdata_pre_5),
	.datad(\D_iw[27]~0_combout ),
	.cin(gnd),
	.combout(\F_iw[5]~21_combout ),
	.cout());
defparam \F_iw[5]~21 .lut_mask = 16'hFEFF;
defparam \F_iw[5]~21 .sum_lutc_input = "datac";

dffeas \D_iw[5] (
	.clk(clk_clk),
	.d(\F_iw[5]~21_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[5]~q ),
	.prn(vcc));
defparam \D_iw[5] .is_wysiwyg = "true";
defparam \D_iw[5] .power_up = "low";

cycloneive_lcell_comb \F_iw[4]~22 (
	.dataa(src_payload6),
	.datab(src1_valid),
	.datac(av_readdata_pre_4),
	.datad(\D_iw[27]~0_combout ),
	.cin(gnd),
	.combout(\F_iw[4]~22_combout ),
	.cout());
defparam \F_iw[4]~22 .lut_mask = 16'hFEFF;
defparam \F_iw[4]~22 .sum_lutc_input = "datac";

dffeas \D_iw[4] (
	.clk(clk_clk),
	.d(\F_iw[4]~22_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[4]~q ),
	.prn(vcc));
defparam \D_iw[4] .is_wysiwyg = "true";
defparam \D_iw[4] .power_up = "low";

cycloneive_lcell_comb \Equal0~7 (
	.dataa(\Equal0~2_combout ),
	.datab(\D_iw[5]~q ),
	.datac(\D_iw[4]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal0~7_combout ),
	.cout());
defparam \Equal0~7 .lut_mask = 16'hFEFE;
defparam \Equal0~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[15]~25 (
	.dataa(src_payload7),
	.datab(src1_valid),
	.datac(av_readdata_pre_15),
	.datad(\D_iw[27]~0_combout ),
	.cin(gnd),
	.combout(\F_iw[15]~25_combout ),
	.cout());
defparam \F_iw[15]~25 .lut_mask = 16'hFEFF;
defparam \F_iw[15]~25 .sum_lutc_input = "datac";

dffeas \D_iw[15] (
	.clk(clk_clk),
	.d(\F_iw[15]~25_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[15]~q ),
	.prn(vcc));
defparam \D_iw[15] .is_wysiwyg = "true";
defparam \D_iw[15] .power_up = "low";

cycloneive_lcell_comb \F_iw[14]~23 (
	.dataa(src1_valid),
	.datab(read_latency_shift_reg_05),
	.datac(q_a_14),
	.datad(av_readdata_pre_14),
	.cin(gnd),
	.combout(\F_iw[14]~23_combout ),
	.cout());
defparam \F_iw[14]~23 .lut_mask = 16'hFFFE;
defparam \F_iw[14]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[14]~24 (
	.dataa(\F_iw[14]~23_combout ),
	.datab(hbreak_enabled1),
	.datac(\hbreak_req~0_combout ),
	.datad(\D_iw[27]~0_combout ),
	.cin(gnd),
	.combout(\F_iw[14]~24_combout ),
	.cout());
defparam \F_iw[14]~24 .lut_mask = 16'hAFCF;
defparam \F_iw[14]~24 .sum_lutc_input = "datac";

dffeas \D_iw[14] (
	.clk(clk_clk),
	.d(\F_iw[14]~24_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[14]~q ),
	.prn(vcc));
defparam \D_iw[14] .is_wysiwyg = "true";
defparam \D_iw[14] .power_up = "low";

cycloneive_lcell_comb \D_op_opx_rsv63~0 (
	.dataa(\D_iw[15]~q ),
	.datab(\D_iw[14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_op_opx_rsv63~0_combout ),
	.cout());
defparam \D_op_opx_rsv63~0 .lut_mask = 16'hEEEE;
defparam \D_op_opx_rsv63~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[13]~11 (
	.dataa(src_payload1),
	.datab(src1_valid),
	.datac(av_readdata_pre_13),
	.datad(\D_iw[27]~0_combout ),
	.cin(gnd),
	.combout(\F_iw[13]~11_combout ),
	.cout());
defparam \F_iw[13]~11 .lut_mask = 16'hFEFF;
defparam \F_iw[13]~11 .sum_lutc_input = "datac";

dffeas \D_iw[13] (
	.clk(clk_clk),
	.d(\F_iw[13]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[13]~q ),
	.prn(vcc));
defparam \D_iw[13] .is_wysiwyg = "true";
defparam \D_iw[13] .power_up = "low";

cycloneive_lcell_comb \F_iw[16]~12 (
	.dataa(src_payload2),
	.datab(src1_valid),
	.datac(av_readdata_pre_16),
	.datad(\D_iw[27]~0_combout ),
	.cin(gnd),
	.combout(\F_iw[16]~12_combout ),
	.cout());
defparam \F_iw[16]~12 .lut_mask = 16'hFEFF;
defparam \F_iw[16]~12 .sum_lutc_input = "datac";

dffeas \D_iw[16] (
	.clk(clk_clk),
	.d(\F_iw[16]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[16]~q ),
	.prn(vcc));
defparam \D_iw[16] .is_wysiwyg = "true";
defparam \D_iw[16] .power_up = "low";

cycloneive_lcell_comb \F_iw[12]~13 (
	.dataa(read_latency_shift_reg_01),
	.datab(mem_73_0),
	.datac(mem_55_0),
	.datad(av_readdata_pre_12),
	.cin(gnd),
	.combout(\F_iw[12]~13_combout ),
	.cout());
defparam \F_iw[12]~13 .lut_mask = 16'hFFFE;
defparam \F_iw[12]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[12]~14 (
	.dataa(\D_iw[27]~0_combout ),
	.datab(\F_iw[12]~13_combout ),
	.datac(read_latency_shift_reg_05),
	.datad(q_a_12),
	.cin(gnd),
	.combout(\F_iw[12]~14_combout ),
	.cout());
defparam \F_iw[12]~14 .lut_mask = 16'hFFFE;
defparam \F_iw[12]~14 .sum_lutc_input = "datac";

dffeas \D_iw[12] (
	.clk(clk_clk),
	.d(\F_iw[12]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[12]~q ),
	.prn(vcc));
defparam \D_iw[12] .is_wysiwyg = "true";
defparam \D_iw[12] .power_up = "low";

cycloneive_lcell_comb \Equal62~4 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~4_combout ),
	.cout());
defparam \Equal62~4 .lut_mask = 16'hFF7F;
defparam \Equal62~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~5 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~5_combout ),
	.cout());
defparam \Equal62~5 .lut_mask = 16'hFFF7;
defparam \Equal62~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~6 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~6_combout ),
	.cout());
defparam \Equal62~6 .lut_mask = 16'hFFFB;
defparam \Equal62~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_shift_rot~0 (
	.dataa(\D_op_opx_rsv63~0_combout ),
	.datab(\Equal62~4_combout ),
	.datac(\Equal62~5_combout ),
	.datad(\Equal62~6_combout ),
	.cin(gnd),
	.combout(\D_ctrl_shift_rot~0_combout ),
	.cout());
defparam \D_ctrl_shift_rot~0 .lut_mask = 16'hFFFE;
defparam \D_ctrl_shift_rot~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_shift_logical~0 (
	.dataa(\D_iw[12]~q ),
	.datab(gnd),
	.datac(\D_iw[13]~q ),
	.datad(\D_iw[16]~q ),
	.cin(gnd),
	.combout(\D_ctrl_shift_logical~0_combout ),
	.cout());
defparam \D_ctrl_shift_logical~0 .lut_mask = 16'hAFFF;
defparam \D_ctrl_shift_logical~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_shift_rot~1 (
	.dataa(\D_ctrl_shift_logical~0_combout ),
	.datab(\Equal62~4_combout ),
	.datac(\D_iw[15]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_ctrl_shift_rot~1_combout ),
	.cout());
defparam \D_ctrl_shift_rot~1 .lut_mask = 16'hACFF;
defparam \D_ctrl_shift_rot~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~7 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~7_combout ),
	.cout());
defparam \Equal62~7 .lut_mask = 16'hFFBF;
defparam \Equal62~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_shift_rot~2 (
	.dataa(\D_ctrl_shift_rot~1_combout ),
	.datab(\Equal62~7_combout ),
	.datac(\D_iw[14]~q ),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_ctrl_shift_rot~2_combout ),
	.cout());
defparam \D_ctrl_shift_rot~2 .lut_mask = 16'hFEFF;
defparam \D_ctrl_shift_rot~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_shift_rot~3 (
	.dataa(\Equal0~7_combout ),
	.datab(\D_ctrl_shift_rot~0_combout ),
	.datac(\D_ctrl_shift_rot~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_shift_rot~3_combout ),
	.cout());
defparam \D_ctrl_shift_rot~3 .lut_mask = 16'hFEFE;
defparam \D_ctrl_shift_rot~3 .sum_lutc_input = "datac";

dffeas R_ctrl_shift_rot(
	.clk(clk_clk),
	.d(\D_ctrl_shift_rot~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_shift_rot~q ),
	.prn(vcc));
defparam R_ctrl_shift_rot.is_wysiwyg = "true";
defparam R_ctrl_shift_rot.power_up = "low";

cycloneive_lcell_comb \E_stall~0 (
	.dataa(\R_ctrl_shift_rot~q ),
	.datab(\E_valid_from_R~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\E_stall~0_combout ),
	.cout());
defparam \E_stall~0 .lut_mask = 16'hEEEE;
defparam \E_stall~0 .sum_lutc_input = "datac";

dffeas E_new_inst(
	.clk(clk_clk),
	.d(\R_valid~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_new_inst~q ),
	.prn(vcc));
defparam E_new_inst.is_wysiwyg = "true";
defparam E_new_inst.power_up = "low";

cycloneive_lcell_comb \E_shift_rot_cnt[0]~5 (
	.dataa(\E_shift_rot_cnt[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\E_shift_rot_cnt[0]~5_combout ),
	.cout(\E_shift_rot_cnt[0]~6 ));
defparam \E_shift_rot_cnt[0]~5 .lut_mask = 16'h55AA;
defparam \E_shift_rot_cnt[0]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_hi_imm16~0 (
	.dataa(\D_iw[0]~q ),
	.datab(\D_iw[1]~q ),
	.datac(\D_iw[4]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\D_ctrl_hi_imm16~0_combout ),
	.cout());
defparam \D_ctrl_hi_imm16~0 .lut_mask = 16'hFFF7;
defparam \D_ctrl_hi_imm16~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_hi_imm16~1 (
	.dataa(\D_iw[2]~q ),
	.datab(\D_iw[5]~q ),
	.datac(\D_ctrl_hi_imm16~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_hi_imm16~1_combout ),
	.cout());
defparam \D_ctrl_hi_imm16~1 .lut_mask = 16'hFEFE;
defparam \D_ctrl_hi_imm16~1 .sum_lutc_input = "datac";

dffeas R_ctrl_hi_imm16(
	.clk(clk_clk),
	.d(\D_ctrl_hi_imm16~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_hi_imm16~q ),
	.prn(vcc));
defparam R_ctrl_hi_imm16.is_wysiwyg = "true";
defparam R_ctrl_hi_imm16.power_up = "low";

cycloneive_lcell_comb \D_ctrl_alu_force_xor~14 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[2]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[0]~q ),
	.cin(gnd),
	.combout(\D_ctrl_alu_force_xor~14_combout ),
	.cout());
defparam \D_ctrl_alu_force_xor~14 .lut_mask = 16'hF6FF;
defparam \D_ctrl_alu_force_xor~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~17 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~17_combout ),
	.cout());
defparam \Equal0~17 .lut_mask = 16'hFFFE;
defparam \Equal0~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~11 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~11_combout ),
	.cout());
defparam \Equal0~11 .lut_mask = 16'hFFFD;
defparam \Equal0~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_force_src2_zero~0 (
	.dataa(\D_iw[5]~q ),
	.datab(\D_ctrl_alu_force_xor~14_combout ),
	.datac(\Equal0~17_combout ),
	.datad(\Equal0~11_combout ),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~0_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~0 .lut_mask = 16'h7FFF;
defparam \D_ctrl_force_src2_zero~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~14 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~14_combout ),
	.cout());
defparam \Equal62~14 .lut_mask = 16'hFEFF;
defparam \Equal62~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~13 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~13_combout ),
	.cout());
defparam \Equal62~13 .lut_mask = 16'hFDFF;
defparam \Equal62~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_force_src2_zero~1 (
	.dataa(\D_iw[15]~q ),
	.datab(\Equal62~14_combout ),
	.datac(\Equal62~13_combout ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~1_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~1 .lut_mask = 16'hFEFF;
defparam \D_ctrl_force_src2_zero~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~11 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~11_combout ),
	.cout());
defparam \Equal62~11 .lut_mask = 16'hEFFF;
defparam \Equal62~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_force_src2_zero~2 (
	.dataa(\Equal0~7_combout ),
	.datab(\D_ctrl_force_src2_zero~1_combout ),
	.datac(\Equal62~11_combout ),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~2_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~2 .lut_mask = 16'hFEFF;
defparam \D_ctrl_force_src2_zero~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~9 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~9_combout ),
	.cout());
defparam \Equal62~9 .lut_mask = 16'hBFFF;
defparam \Equal62~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_force_src2_zero~3 (
	.dataa(\D_iw[15]~q ),
	.datab(gnd),
	.datac(\Equal0~7_combout ),
	.datad(\Equal62~9_combout ),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~3_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~3 .lut_mask = 16'hAFFF;
defparam \D_ctrl_force_src2_zero~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~12 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~12_combout ),
	.cout());
defparam \Equal0~12 .lut_mask = 16'hDFFF;
defparam \Equal0~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~8 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~8_combout ),
	.cout());
defparam \Equal62~8 .lut_mask = 16'hFFEF;
defparam \Equal62~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~3 (
	.dataa(\D_iw[5]~q ),
	.datab(\D_iw[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal0~3_combout ),
	.cout());
defparam \Equal0~3 .lut_mask = 16'hEEEE;
defparam \Equal0~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_op_cmpge~0 (
	.dataa(\Equal0~2_combout ),
	.datab(\Equal0~3_combout ),
	.datac(\D_iw[14]~q ),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_op_cmpge~0_combout ),
	.cout());
defparam \D_op_cmpge~0 .lut_mask = 16'hFEFF;
defparam \D_op_cmpge~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_implicit_dst_eretaddr~1 (
	.dataa(gnd),
	.datab(\Equal62~4_combout ),
	.datac(\Equal62~8_combout ),
	.datad(\D_op_cmpge~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~1_combout ),
	.cout());
defparam \D_ctrl_implicit_dst_eretaddr~1 .lut_mask = 16'h3FFF;
defparam \D_ctrl_implicit_dst_eretaddr~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~10 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~10_combout ),
	.cout());
defparam \Equal62~10 .lut_mask = 16'hDFFF;
defparam \Equal62~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_op_opx_rsv17~0 (
	.dataa(\Equal0~2_combout ),
	.datab(\Equal0~3_combout ),
	.datac(\D_iw[15]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_op_opx_rsv17~0_combout ),
	.cout());
defparam \D_op_opx_rsv17~0 .lut_mask = 16'hFEFF;
defparam \D_op_opx_rsv17~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_implicit_dst_eretaddr~2 (
	.dataa(gnd),
	.datab(\Equal62~9_combout ),
	.datac(\Equal62~10_combout ),
	.datad(\D_op_opx_rsv17~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~2_combout ),
	.cout());
defparam \D_ctrl_implicit_dst_eretaddr~2 .lut_mask = 16'h3FFF;
defparam \D_ctrl_implicit_dst_eretaddr~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~2 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~2_combout ),
	.cout());
defparam \Equal62~2 .lut_mask = 16'hFBFF;
defparam \Equal62~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_op_opx_rsv00~0 (
	.dataa(\Equal0~2_combout ),
	.datab(\Equal0~3_combout ),
	.datac(\D_iw[15]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_op_opx_rsv00~0_combout ),
	.cout());
defparam \D_op_opx_rsv00~0 .lut_mask = 16'hEFFF;
defparam \D_op_opx_rsv00~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_implicit_dst_eretaddr~3 (
	.dataa(gnd),
	.datab(\Equal62~2_combout ),
	.datac(\Equal62~0_combout ),
	.datad(\D_op_opx_rsv00~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~3_combout ),
	.cout());
defparam \D_ctrl_implicit_dst_eretaddr~3 .lut_mask = 16'h3FFF;
defparam \D_ctrl_implicit_dst_eretaddr~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_implicit_dst_eretaddr~4 (
	.dataa(gnd),
	.datab(\Equal62~5_combout ),
	.datac(\Equal62~6_combout ),
	.datad(\D_op_opx_rsv00~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~4_combout ),
	.cout());
defparam \D_ctrl_implicit_dst_eretaddr~4 .lut_mask = 16'h3FFF;
defparam \D_ctrl_implicit_dst_eretaddr~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_implicit_dst_eretaddr~5 (
	.dataa(\D_ctrl_implicit_dst_eretaddr~1_combout ),
	.datab(\D_ctrl_implicit_dst_eretaddr~2_combout ),
	.datac(\D_ctrl_implicit_dst_eretaddr~3_combout ),
	.datad(\D_ctrl_implicit_dst_eretaddr~4_combout ),
	.cin(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~5_combout ),
	.cout());
defparam \D_ctrl_implicit_dst_eretaddr~5 .lut_mask = 16'hFFFE;
defparam \D_ctrl_implicit_dst_eretaddr~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_implicit_dst_eretaddr~6 (
	.dataa(\Equal62~5_combout ),
	.datab(\Equal62~11_combout ),
	.datac(\D_op_opx_rsv17~0_combout ),
	.datad(\D_op_cmpge~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~6_combout ),
	.cout());
defparam \D_ctrl_implicit_dst_eretaddr~6 .lut_mask = 16'h7FFF;
defparam \D_ctrl_implicit_dst_eretaddr~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~1 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~1_combout ),
	.cout());
defparam \Equal62~1 .lut_mask = 16'hF7FF;
defparam \Equal62~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~12 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~12_combout ),
	.cout());
defparam \Equal62~12 .lut_mask = 16'hFFFE;
defparam \Equal62~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_implicit_dst_eretaddr~7 (
	.dataa(\D_iw[15]~q ),
	.datab(\D_iw[14]~q ),
	.datac(\Equal62~12_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~7_combout ),
	.cout());
defparam \D_ctrl_implicit_dst_eretaddr~7 .lut_mask = 16'h7F7F;
defparam \D_ctrl_implicit_dst_eretaddr~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_implicit_dst_eretaddr~8 (
	.dataa(\Equal62~1_combout ),
	.datab(\Equal62~9_combout ),
	.datac(\D_op_opx_rsv63~0_combout ),
	.datad(\D_ctrl_implicit_dst_eretaddr~7_combout ),
	.cin(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~8_combout ),
	.cout());
defparam \D_ctrl_implicit_dst_eretaddr~8 .lut_mask = 16'hFF7F;
defparam \D_ctrl_implicit_dst_eretaddr~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_implicit_dst_eretaddr~9 (
	.dataa(\Equal62~6_combout ),
	.datab(\D_op_cmpge~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~9_combout ),
	.cout());
defparam \D_ctrl_implicit_dst_eretaddr~9 .lut_mask = 16'h7777;
defparam \D_ctrl_implicit_dst_eretaddr~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_implicit_dst_eretaddr~10 (
	.dataa(\Equal0~7_combout ),
	.datab(\D_ctrl_implicit_dst_eretaddr~6_combout ),
	.datac(\D_ctrl_implicit_dst_eretaddr~8_combout ),
	.datad(\D_ctrl_implicit_dst_eretaddr~9_combout ),
	.cin(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~10_combout ),
	.cout());
defparam \D_ctrl_implicit_dst_eretaddr~10 .lut_mask = 16'hFFFD;
defparam \D_ctrl_implicit_dst_eretaddr~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal62~3 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~3_combout ),
	.cout());
defparam \Equal62~3 .lut_mask = 16'hFFFD;
defparam \Equal62~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_implicit_dst_eretaddr~11 (
	.dataa(\Equal62~3_combout ),
	.datab(\Equal62~13_combout ),
	.datac(\Equal0~7_combout ),
	.datad(\D_op_opx_rsv63~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~11_combout ),
	.cout());
defparam \D_ctrl_implicit_dst_eretaddr~11 .lut_mask = 16'h7FFF;
defparam \D_ctrl_implicit_dst_eretaddr~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~15 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~15_combout ),
	.cout());
defparam \Equal0~15 .lut_mask = 16'hFDFF;
defparam \Equal0~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_implicit_dst_eretaddr~12 (
	.dataa(\D_ctrl_implicit_dst_eretaddr~11_combout ),
	.datab(\Equal62~6_combout ),
	.datac(\D_op_opx_rsv17~0_combout ),
	.datad(\Equal0~15_combout ),
	.cin(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~12_combout ),
	.cout());
defparam \D_ctrl_implicit_dst_eretaddr~12 .lut_mask = 16'hBFFF;
defparam \D_ctrl_implicit_dst_eretaddr~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~4 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~4_combout ),
	.cout());
defparam \Equal0~4 .lut_mask = 16'h7FFF;
defparam \Equal0~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~16 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~16_combout ),
	.cout());
defparam \Equal0~16 .lut_mask = 16'hBFFF;
defparam \Equal0~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_force_src2_zero~4 (
	.dataa(\D_iw[5]~q ),
	.datab(\D_iw[4]~q ),
	.datac(\Equal0~4_combout ),
	.datad(\Equal0~16_combout ),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~4_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~4 .lut_mask = 16'hEFFF;
defparam \D_ctrl_force_src2_zero~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_retaddr~0 (
	.dataa(\D_iw[15]~q ),
	.datab(\Equal62~10_combout ),
	.datac(\Equal62~11_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~0_combout ),
	.cout());
defparam \D_ctrl_retaddr~0 .lut_mask = 16'hFEFE;
defparam \D_ctrl_retaddr~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_retaddr~1 (
	.dataa(\Equal62~13_combout ),
	.datab(\Equal62~14_combout ),
	.datac(gnd),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~1_combout ),
	.cout());
defparam \D_ctrl_retaddr~1 .lut_mask = 16'hEEFF;
defparam \D_ctrl_retaddr~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_retaddr~2 (
	.dataa(\Equal0~7_combout ),
	.datab(\D_iw[14]~q ),
	.datac(\D_ctrl_retaddr~0_combout ),
	.datad(\D_ctrl_retaddr~1_combout ),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~2_combout ),
	.cout());
defparam \D_ctrl_retaddr~2 .lut_mask = 16'hFFFE;
defparam \D_ctrl_retaddr~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_force_src2_zero~5 (
	.dataa(\D_ctrl_force_src2_zero~4_combout ),
	.datab(\D_iw[5]~q ),
	.datac(\Equal0~2_combout ),
	.datad(\D_ctrl_retaddr~2_combout ),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~5_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~5 .lut_mask = 16'hEFFF;
defparam \D_ctrl_force_src2_zero~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_force_src2_zero~6 (
	.dataa(\D_ctrl_implicit_dst_eretaddr~5_combout ),
	.datab(\D_ctrl_implicit_dst_eretaddr~10_combout ),
	.datac(\D_ctrl_implicit_dst_eretaddr~12_combout ),
	.datad(\D_ctrl_force_src2_zero~5_combout ),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~6_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~6 .lut_mask = 16'hFFFE;
defparam \D_ctrl_force_src2_zero~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_force_src2_zero~7 (
	.dataa(\D_ctrl_force_src2_zero~2_combout ),
	.datab(\D_ctrl_force_src2_zero~3_combout ),
	.datac(\Equal0~12_combout ),
	.datad(\D_ctrl_force_src2_zero~6_combout ),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~7_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~7 .lut_mask = 16'hFFDF;
defparam \D_ctrl_force_src2_zero~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_force_src2_zero~8 (
	.dataa(\D_iw[4]~q ),
	.datab(\Equal0~16_combout ),
	.datac(\D_iw[5]~q ),
	.datad(\Equal0~2_combout ),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~8_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~8 .lut_mask = 16'hFFDE;
defparam \D_ctrl_force_src2_zero~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_force_src2_zero~9 (
	.dataa(\D_ctrl_force_src2_zero~0_combout ),
	.datab(\D_ctrl_force_src2_zero~7_combout ),
	.datac(\D_iw[4]~q ),
	.datad(\D_ctrl_force_src2_zero~8_combout ),
	.cin(gnd),
	.combout(\D_ctrl_force_src2_zero~9_combout ),
	.cout());
defparam \D_ctrl_force_src2_zero~9 .lut_mask = 16'hFFF7;
defparam \D_ctrl_force_src2_zero~9 .sum_lutc_input = "datac";

dffeas R_ctrl_force_src2_zero(
	.clk(clk_clk),
	.d(\D_ctrl_force_src2_zero~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_force_src2_zero~q ),
	.prn(vcc));
defparam R_ctrl_force_src2_zero.is_wysiwyg = "true";
defparam R_ctrl_force_src2_zero.power_up = "low";

cycloneive_lcell_comb \R_src2_lo[3]~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\R_ctrl_hi_imm16~q ),
	.datad(\R_ctrl_force_src2_zero~q ),
	.cin(gnd),
	.combout(\R_src2_lo[3]~8_combout ),
	.cout());
defparam \R_src2_lo[3]~8 .lut_mask = 16'h0FFF;
defparam \R_src2_lo[3]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[6]~38 (
	.dataa(read_latency_shift_reg_01),
	.datab(mem_73_0),
	.datac(mem_55_0),
	.datad(av_readdata_pre_6),
	.cin(gnd),
	.combout(\F_iw[6]~38_combout ),
	.cout());
defparam \F_iw[6]~38 .lut_mask = 16'hFFFE;
defparam \F_iw[6]~38 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[6]~39 (
	.dataa(\D_iw[27]~0_combout ),
	.datab(\F_iw[6]~38_combout ),
	.datac(read_latency_shift_reg_05),
	.datad(q_a_6),
	.cin(gnd),
	.combout(\F_iw[6]~39_combout ),
	.cout());
defparam \F_iw[6]~39 .lut_mask = 16'hFFFE;
defparam \F_iw[6]~39 .sum_lutc_input = "datac";

dffeas \D_iw[6] (
	.clk(clk_clk),
	.d(\F_iw[6]~39_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[6]~q ),
	.prn(vcc));
defparam \D_iw[6] .is_wysiwyg = "true";
defparam \D_iw[6] .power_up = "low";

cycloneive_lcell_comb \D_ctrl_implicit_dst_eretaddr~0 (
	.dataa(\D_iw[14]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~0_combout ),
	.cout());
defparam \D_ctrl_implicit_dst_eretaddr~0 .lut_mask = 16'hAAFF;
defparam \D_ctrl_implicit_dst_eretaddr~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_unsigned_lo_imm16~2 (
	.dataa(\D_op_opx_rsv63~0_combout ),
	.datab(\Equal62~5_combout ),
	.datac(\Equal62~4_combout ),
	.datad(\D_ctrl_implicit_dst_eretaddr~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_unsigned_lo_imm16~2_combout ),
	.cout());
defparam \D_ctrl_unsigned_lo_imm16~2 .lut_mask = 16'hFEFF;
defparam \D_ctrl_unsigned_lo_imm16~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_unsigned_lo_imm16~5 (
	.dataa(\Equal0~2_combout ),
	.datab(\D_iw[5]~q ),
	.datac(\D_iw[4]~q ),
	.datad(\D_ctrl_unsigned_lo_imm16~2_combout ),
	.cin(gnd),
	.combout(\D_ctrl_unsigned_lo_imm16~5_combout ),
	.cout());
defparam \D_ctrl_unsigned_lo_imm16~5 .lut_mask = 16'hFFFE;
defparam \D_ctrl_unsigned_lo_imm16~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_b_is_dst~0 (
	.dataa(\D_iw[2]~q ),
	.datab(\D_iw[3]~q ),
	.datac(\D_iw[5]~q ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_b_is_dst~0_combout ),
	.cout());
defparam \D_ctrl_b_is_dst~0 .lut_mask = 16'h6996;
defparam \D_ctrl_b_is_dst~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_b_is_dst~1 (
	.dataa(\D_iw[2]~q ),
	.datab(\D_iw[3]~q ),
	.datac(\D_iw[5]~q ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_b_is_dst~1_combout ),
	.cout());
defparam \D_ctrl_b_is_dst~1 .lut_mask = 16'hFBFE;
defparam \D_ctrl_b_is_dst~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_b_is_dst~2 (
	.dataa(\D_iw[0]~q ),
	.datab(\D_iw[1]~q ),
	.datac(\D_ctrl_b_is_dst~0_combout ),
	.datad(\D_ctrl_b_is_dst~1_combout ),
	.cin(gnd),
	.combout(\D_ctrl_b_is_dst~2_combout ),
	.cout());
defparam \D_ctrl_b_is_dst~2 .lut_mask = 16'h96FF;
defparam \D_ctrl_b_is_dst~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~13 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~13_combout ),
	.cout());
defparam \Equal0~13 .lut_mask = 16'hFFDF;
defparam \Equal0~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_use_imm~0 (
	.dataa(\D_ctrl_b_is_dst~2_combout ),
	.datab(\Equal0~13_combout ),
	.datac(\Equal0~11_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\R_src2_use_imm~0_combout ),
	.cout());
defparam \R_src2_use_imm~0 .lut_mask = 16'hFEFF;
defparam \R_src2_use_imm~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_ctrl_br_nxt~0 (
	.dataa(\D_iw[0]~q ),
	.datab(\D_iw[4]~q ),
	.datac(\D_iw[5]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\R_ctrl_br_nxt~0_combout ),
	.cout());
defparam \R_ctrl_br_nxt~0 .lut_mask = 16'hFFFE;
defparam \R_ctrl_br_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_ctrl_br_nxt~1 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[2]~q ),
	.datac(gnd),
	.datad(\R_ctrl_br_nxt~0_combout ),
	.cin(gnd),
	.combout(\R_ctrl_br_nxt~1_combout ),
	.cout());
defparam \R_ctrl_br_nxt~1 .lut_mask = 16'hEEFF;
defparam \R_ctrl_br_nxt~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_use_imm~1 (
	.dataa(\D_ctrl_unsigned_lo_imm16~5_combout ),
	.datab(\R_src2_use_imm~0_combout ),
	.datac(\R_valid~q ),
	.datad(\R_ctrl_br_nxt~1_combout ),
	.cin(gnd),
	.combout(\R_src2_use_imm~1_combout ),
	.cout());
defparam \R_src2_use_imm~1 .lut_mask = 16'hFFFE;
defparam \R_src2_use_imm~1 .sum_lutc_input = "datac";

dffeas R_src2_use_imm(
	.clk(clk_clk),
	.d(\R_src2_use_imm~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_src2_use_imm~q ),
	.prn(vcc));
defparam R_src2_use_imm.is_wysiwyg = "true";
defparam R_src2_use_imm.power_up = "low";

cycloneive_lcell_comb \D_ctrl_src_imm5_shift_rot~0 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[15]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_ctrl_src_imm5_shift_rot~0_combout ),
	.cout());
defparam \D_ctrl_src_imm5_shift_rot~0 .lut_mask = 16'hBBF3;
defparam \D_ctrl_src_imm5_shift_rot~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_src_imm5_shift_rot~1 (
	.dataa(\Equal0~7_combout ),
	.datab(\D_iw[12]~q ),
	.datac(\D_iw[13]~q ),
	.datad(\D_ctrl_src_imm5_shift_rot~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_src_imm5_shift_rot~1_combout ),
	.cout());
defparam \D_ctrl_src_imm5_shift_rot~1 .lut_mask = 16'hEFFF;
defparam \D_ctrl_src_imm5_shift_rot~1 .sum_lutc_input = "datac";

dffeas R_ctrl_src_imm5_shift_rot(
	.clk(clk_clk),
	.d(\D_ctrl_src_imm5_shift_rot~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_src_imm5_shift_rot~q ),
	.prn(vcc));
defparam R_ctrl_src_imm5_shift_rot.is_wysiwyg = "true";
defparam R_ctrl_src_imm5_shift_rot.power_up = "low";

cycloneive_lcell_comb \R_src2_lo~9 (
	.dataa(\R_src2_use_imm~q ),
	.datab(\R_ctrl_src_imm5_shift_rot~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\R_src2_lo~9_combout ),
	.cout());
defparam \R_src2_lo~9 .lut_mask = 16'hEEEE;
defparam \R_src2_lo~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_lo[0]~14 (
	.dataa(\R_src2_lo[3]~8_combout ),
	.datab(\D_iw[6]~q ),
	.datac(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.datad(\R_src2_lo~9_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[0]~14_combout ),
	.cout());
defparam \R_src2_lo[0]~14 .lut_mask = 16'hFAFC;
defparam \R_src2_lo[0]~14 .sum_lutc_input = "datac";

dffeas \E_src2[0] (
	.clk(clk_clk),
	.d(\R_src2_lo[0]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[0]~q ),
	.prn(vcc));
defparam \E_src2[0] .is_wysiwyg = "true";
defparam \E_src2[0] .power_up = "low";

dffeas \E_shift_rot_cnt[0] (
	.clk(clk_clk),
	.d(\E_shift_rot_cnt[0]~5_combout ),
	.asdata(\E_src2[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_cnt[0]~q ),
	.prn(vcc));
defparam \E_shift_rot_cnt[0] .is_wysiwyg = "true";
defparam \E_shift_rot_cnt[0] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_cnt[1]~7 (
	.dataa(\E_shift_rot_cnt[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\E_shift_rot_cnt[0]~6 ),
	.combout(\E_shift_rot_cnt[1]~7_combout ),
	.cout(\E_shift_rot_cnt[1]~8 ));
defparam \E_shift_rot_cnt[1]~7 .lut_mask = 16'h5A5F;
defparam \E_shift_rot_cnt[1]~7 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_iw[7]~36 (
	.dataa(read_latency_shift_reg_01),
	.datab(mem_73_0),
	.datac(mem_55_0),
	.datad(av_readdata_pre_7),
	.cin(gnd),
	.combout(\F_iw[7]~36_combout ),
	.cout());
defparam \F_iw[7]~36 .lut_mask = 16'hFFFE;
defparam \F_iw[7]~36 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[7]~37 (
	.dataa(\D_iw[27]~0_combout ),
	.datab(\F_iw[7]~36_combout ),
	.datac(read_latency_shift_reg_05),
	.datad(q_a_7),
	.cin(gnd),
	.combout(\F_iw[7]~37_combout ),
	.cout());
defparam \F_iw[7]~37 .lut_mask = 16'hFFFE;
defparam \F_iw[7]~37 .sum_lutc_input = "datac";

dffeas \D_iw[7] (
	.clk(clk_clk),
	.d(\F_iw[7]~37_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[7]~q ),
	.prn(vcc));
defparam \D_iw[7] .is_wysiwyg = "true";
defparam \D_iw[7] .power_up = "low";

cycloneive_lcell_comb \R_src2_lo[1]~13 (
	.dataa(\R_src2_lo[3]~8_combout ),
	.datab(\D_iw[7]~q ),
	.datac(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.datad(\R_src2_lo~9_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[1]~13_combout ),
	.cout());
defparam \R_src2_lo[1]~13 .lut_mask = 16'hFAFC;
defparam \R_src2_lo[1]~13 .sum_lutc_input = "datac";

dffeas \E_src2[1] (
	.clk(clk_clk),
	.d(\R_src2_lo[1]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[1]~q ),
	.prn(vcc));
defparam \E_src2[1] .is_wysiwyg = "true";
defparam \E_src2[1] .power_up = "low";

dffeas \E_shift_rot_cnt[1] (
	.clk(clk_clk),
	.d(\E_shift_rot_cnt[1]~7_combout ),
	.asdata(\E_src2[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_cnt[1]~q ),
	.prn(vcc));
defparam \E_shift_rot_cnt[1] .is_wysiwyg = "true";
defparam \E_shift_rot_cnt[1] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_cnt[2]~9 (
	.dataa(\E_shift_rot_cnt[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\E_shift_rot_cnt[1]~8 ),
	.combout(\E_shift_rot_cnt[2]~9_combout ),
	.cout(\E_shift_rot_cnt[2]~10 ));
defparam \E_shift_rot_cnt[2]~9 .lut_mask = 16'h5AAF;
defparam \E_shift_rot_cnt[2]~9 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_iw[8]~34 (
	.dataa(read_latency_shift_reg_01),
	.datab(mem_73_0),
	.datac(mem_55_0),
	.datad(av_readdata_pre_8),
	.cin(gnd),
	.combout(\F_iw[8]~34_combout ),
	.cout());
defparam \F_iw[8]~34 .lut_mask = 16'hFFFE;
defparam \F_iw[8]~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[8]~35 (
	.dataa(\D_iw[27]~0_combout ),
	.datab(\F_iw[8]~34_combout ),
	.datac(read_latency_shift_reg_05),
	.datad(q_a_8),
	.cin(gnd),
	.combout(\F_iw[8]~35_combout ),
	.cout());
defparam \F_iw[8]~35 .lut_mask = 16'hFFFE;
defparam \F_iw[8]~35 .sum_lutc_input = "datac";

dffeas \D_iw[8] (
	.clk(clk_clk),
	.d(\F_iw[8]~35_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[8]~q ),
	.prn(vcc));
defparam \D_iw[8] .is_wysiwyg = "true";
defparam \D_iw[8] .power_up = "low";

cycloneive_lcell_comb \R_src2_lo[2]~12 (
	.dataa(\R_src2_lo[3]~8_combout ),
	.datab(\D_iw[8]~q ),
	.datac(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.datad(\R_src2_lo~9_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[2]~12_combout ),
	.cout());
defparam \R_src2_lo[2]~12 .lut_mask = 16'hFAFC;
defparam \R_src2_lo[2]~12 .sum_lutc_input = "datac";

dffeas \E_src2[2] (
	.clk(clk_clk),
	.d(\R_src2_lo[2]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[2]~q ),
	.prn(vcc));
defparam \E_src2[2] .is_wysiwyg = "true";
defparam \E_src2[2] .power_up = "low";

dffeas \E_shift_rot_cnt[2] (
	.clk(clk_clk),
	.d(\E_shift_rot_cnt[2]~9_combout ),
	.asdata(\E_src2[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_cnt[2]~q ),
	.prn(vcc));
defparam \E_shift_rot_cnt[2] .is_wysiwyg = "true";
defparam \E_shift_rot_cnt[2] .power_up = "low";

cycloneive_lcell_comb \E_stall~1 (
	.dataa(\E_new_inst~q ),
	.datab(\E_shift_rot_cnt[0]~q ),
	.datac(\E_shift_rot_cnt[1]~q ),
	.datad(\E_shift_rot_cnt[2]~q ),
	.cin(gnd),
	.combout(\E_stall~1_combout ),
	.cout());
defparam \E_stall~1 .lut_mask = 16'hFFFE;
defparam \E_stall~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_shift_rot_cnt[3]~11 (
	.dataa(\E_shift_rot_cnt[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\E_shift_rot_cnt[2]~10 ),
	.combout(\E_shift_rot_cnt[3]~11_combout ),
	.cout(\E_shift_rot_cnt[3]~12 ));
defparam \E_shift_rot_cnt[3]~11 .lut_mask = 16'h5A5F;
defparam \E_shift_rot_cnt[3]~11 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_iw[9]~32 (
	.dataa(read_latency_shift_reg_01),
	.datab(mem_73_0),
	.datac(mem_55_0),
	.datad(av_readdata_pre_9),
	.cin(gnd),
	.combout(\F_iw[9]~32_combout ),
	.cout());
defparam \F_iw[9]~32 .lut_mask = 16'hFFFE;
defparam \F_iw[9]~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[9]~33 (
	.dataa(\D_iw[27]~0_combout ),
	.datab(\F_iw[9]~32_combout ),
	.datac(read_latency_shift_reg_05),
	.datad(q_a_9),
	.cin(gnd),
	.combout(\F_iw[9]~33_combout ),
	.cout());
defparam \F_iw[9]~33 .lut_mask = 16'hFFFE;
defparam \F_iw[9]~33 .sum_lutc_input = "datac";

dffeas \D_iw[9] (
	.clk(clk_clk),
	.d(\F_iw[9]~33_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[9]~q ),
	.prn(vcc));
defparam \D_iw[9] .is_wysiwyg = "true";
defparam \D_iw[9] .power_up = "low";

cycloneive_lcell_comb \R_src2_lo[3]~11 (
	.dataa(\R_src2_lo[3]~8_combout ),
	.datab(\D_iw[9]~q ),
	.datac(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.datad(\R_src2_lo~9_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[3]~11_combout ),
	.cout());
defparam \R_src2_lo[3]~11 .lut_mask = 16'hFAFC;
defparam \R_src2_lo[3]~11 .sum_lutc_input = "datac";

dffeas \E_src2[3] (
	.clk(clk_clk),
	.d(\R_src2_lo[3]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[3]~q ),
	.prn(vcc));
defparam \E_src2[3] .is_wysiwyg = "true";
defparam \E_src2[3] .power_up = "low";

dffeas \E_shift_rot_cnt[3] (
	.clk(clk_clk),
	.d(\E_shift_rot_cnt[3]~11_combout ),
	.asdata(\E_src2[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_cnt[3]~q ),
	.prn(vcc));
defparam \E_shift_rot_cnt[3] .is_wysiwyg = "true";
defparam \E_shift_rot_cnt[3] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_cnt[4]~13 (
	.dataa(\E_shift_rot_cnt[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\E_shift_rot_cnt[3]~12 ),
	.combout(\E_shift_rot_cnt[4]~13_combout ),
	.cout());
defparam \E_shift_rot_cnt[4]~13 .lut_mask = 16'h5A5A;
defparam \E_shift_rot_cnt[4]~13 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_iw[10]~30 (
	.dataa(read_latency_shift_reg_01),
	.datab(mem_73_0),
	.datac(mem_55_0),
	.datad(av_readdata_pre_10),
	.cin(gnd),
	.combout(\F_iw[10]~30_combout ),
	.cout());
defparam \F_iw[10]~30 .lut_mask = 16'hFFFE;
defparam \F_iw[10]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[10]~31 (
	.dataa(\D_iw[27]~0_combout ),
	.datab(\F_iw[10]~30_combout ),
	.datac(read_latency_shift_reg_05),
	.datad(q_a_10),
	.cin(gnd),
	.combout(\F_iw[10]~31_combout ),
	.cout());
defparam \F_iw[10]~31 .lut_mask = 16'hFFFE;
defparam \F_iw[10]~31 .sum_lutc_input = "datac";

dffeas \D_iw[10] (
	.clk(clk_clk),
	.d(\F_iw[10]~31_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[10]~q ),
	.prn(vcc));
defparam \D_iw[10] .is_wysiwyg = "true";
defparam \D_iw[10] .power_up = "low";

cycloneive_lcell_comb \R_src2_lo[4]~10 (
	.dataa(\R_src2_lo[3]~8_combout ),
	.datab(\D_iw[10]~q ),
	.datac(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.datad(\R_src2_lo~9_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[4]~10_combout ),
	.cout());
defparam \R_src2_lo[4]~10 .lut_mask = 16'hFAFC;
defparam \R_src2_lo[4]~10 .sum_lutc_input = "datac";

dffeas \E_src2[4] (
	.clk(clk_clk),
	.d(\R_src2_lo[4]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[4]~q ),
	.prn(vcc));
defparam \E_src2[4] .is_wysiwyg = "true";
defparam \E_src2[4] .power_up = "low";

dffeas \E_shift_rot_cnt[4] (
	.clk(clk_clk),
	.d(\E_shift_rot_cnt[4]~13_combout ),
	.asdata(\E_src2[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_cnt[4]~q ),
	.prn(vcc));
defparam \E_shift_rot_cnt[4] .is_wysiwyg = "true";
defparam \E_shift_rot_cnt[4] .power_up = "low";

cycloneive_lcell_comb \E_stall~2 (
	.dataa(\E_stall~0_combout ),
	.datab(\E_stall~1_combout ),
	.datac(\E_shift_rot_cnt[3]~q ),
	.datad(\E_shift_rot_cnt[4]~q ),
	.cin(gnd),
	.combout(\E_stall~2_combout ),
	.cout());
defparam \E_stall~2 .lut_mask = 16'hFFFE;
defparam \E_stall~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_st~0 (
	.dataa(\D_iw[0]~q ),
	.datab(\D_iw[1]~q ),
	.datac(\D_iw[4]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\D_ctrl_st~0_combout ),
	.cout());
defparam \D_ctrl_st~0 .lut_mask = 16'hBFFF;
defparam \D_ctrl_st~0 .sum_lutc_input = "datac";

dffeas R_ctrl_st(
	.clk(clk_clk),
	.d(\D_ctrl_st~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(!\D_iw[2]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_st~q ),
	.prn(vcc));
defparam R_ctrl_st.is_wysiwyg = "true";
defparam R_ctrl_st.power_up = "low";

cycloneive_lcell_comb \D_ctrl_ld_signed~0 (
	.dataa(\D_iw[0]~q ),
	.datab(\D_iw[1]~q ),
	.datac(\D_iw[4]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\D_ctrl_ld_signed~0_combout ),
	.cout());
defparam \D_ctrl_ld_signed~0 .lut_mask = 16'hEFFF;
defparam \D_ctrl_ld_signed~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_ld~2 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[2]~q ),
	.datac(\D_iw[4]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_ld~2_combout ),
	.cout());
defparam \D_ctrl_ld~2 .lut_mask = 16'hBFBF;
defparam \D_ctrl_ld~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_ld~3 (
	.dataa(\D_iw[2]~q ),
	.datab(\D_ctrl_ld_signed~0_combout ),
	.datac(\D_iw[0]~q ),
	.datad(\D_ctrl_ld~2_combout ),
	.cin(gnd),
	.combout(\D_ctrl_ld~3_combout ),
	.cout());
defparam \D_ctrl_ld~3 .lut_mask = 16'hFFFE;
defparam \D_ctrl_ld~3 .sum_lutc_input = "datac";

dffeas R_ctrl_ld(
	.clk(clk_clk),
	.d(\D_ctrl_ld~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_ld~q ),
	.prn(vcc));
defparam R_ctrl_ld.is_wysiwyg = "true";
defparam R_ctrl_ld.power_up = "low";

dffeas av_ld_waiting_for_data(
	.clk(clk_clk),
	.d(\av_ld_waiting_for_data_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_waiting_for_data~q ),
	.prn(vcc));
defparam av_ld_waiting_for_data.is_wysiwyg = "true";
defparam av_ld_waiting_for_data.power_up = "low";

cycloneive_lcell_comb \av_ld_waiting_for_data_nxt~0 (
	.dataa(\E_new_inst~q ),
	.datab(\R_ctrl_ld~q ),
	.datac(\av_ld_waiting_for_data~q ),
	.datad(d_read1),
	.cin(gnd),
	.combout(\av_ld_waiting_for_data_nxt~0_combout ),
	.cout());
defparam \av_ld_waiting_for_data_nxt~0 .lut_mask = 16'hACFF;
defparam \av_ld_waiting_for_data_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_waiting_for_data_nxt~1 (
	.dataa(\av_ld_waiting_for_data_nxt~0_combout ),
	.datab(WideOr1),
	.datac(WideOr13),
	.datad(\av_ld_waiting_for_data~q ),
	.cin(gnd),
	.combout(\av_ld_waiting_for_data_nxt~1_combout ),
	.cout());
defparam \av_ld_waiting_for_data_nxt~1 .lut_mask = 16'hFFFE;
defparam \av_ld_waiting_for_data_nxt~1 .sum_lutc_input = "datac";

dffeas av_ld_aligning_data(
	.clk(clk_clk),
	.d(\av_ld_aligning_data_nxt~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_aligning_data~q ),
	.prn(vcc));
defparam av_ld_aligning_data.is_wysiwyg = "true";
defparam av_ld_aligning_data.power_up = "low";

cycloneive_lcell_comb \av_ld_align_cycle_nxt[0]~0 (
	.dataa(\av_ld_align_cycle[0]~q ),
	.datab(d_read1),
	.datac(WideOr1),
	.datad(WideOr13),
	.cin(gnd),
	.combout(\av_ld_align_cycle_nxt[0]~0_combout ),
	.cout());
defparam \av_ld_align_cycle_nxt[0]~0 .lut_mask = 16'hFFF7;
defparam \av_ld_align_cycle_nxt[0]~0 .sum_lutc_input = "datac";

dffeas \av_ld_align_cycle[0] (
	.clk(clk_clk),
	.d(\av_ld_align_cycle_nxt[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_align_cycle[0]~q ),
	.prn(vcc));
defparam \av_ld_align_cycle[0] .is_wysiwyg = "true";
defparam \av_ld_align_cycle[0] .power_up = "low";

cycloneive_lcell_comb \D_ctrl_mem16~0 (
	.dataa(\D_iw[0]~q ),
	.datab(\D_iw[1]~q ),
	.datac(\D_iw[2]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\D_ctrl_mem16~0_combout ),
	.cout());
defparam \D_ctrl_mem16~0 .lut_mask = 16'hFFFE;
defparam \D_ctrl_mem16~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_mem16~1 (
	.dataa(\D_ctrl_mem16~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_mem16~1_combout ),
	.cout());
defparam \D_ctrl_mem16~1 .lut_mask = 16'hAAFF;
defparam \D_ctrl_mem16~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_align_cycle_nxt[1]~1 (
	.dataa(WideOr11),
	.datab(d_read1),
	.datac(\av_ld_align_cycle[1]~q ),
	.datad(\av_ld_align_cycle[0]~q ),
	.cin(gnd),
	.combout(\av_ld_align_cycle_nxt[1]~1_combout ),
	.cout());
defparam \av_ld_align_cycle_nxt[1]~1 .lut_mask = 16'hBFFB;
defparam \av_ld_align_cycle_nxt[1]~1 .sum_lutc_input = "datac";

dffeas \av_ld_align_cycle[1] (
	.clk(clk_clk),
	.d(\av_ld_align_cycle_nxt[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_align_cycle[1]~q ),
	.prn(vcc));
defparam \av_ld_align_cycle[1] .is_wysiwyg = "true";
defparam \av_ld_align_cycle[1] .power_up = "low";

cycloneive_lcell_comb \av_ld_aligning_data_nxt~0 (
	.dataa(\av_ld_aligning_data~q ),
	.datab(\av_ld_align_cycle[0]~q ),
	.datac(\D_ctrl_mem16~1_combout ),
	.datad(\av_ld_align_cycle[1]~q ),
	.cin(gnd),
	.combout(\av_ld_aligning_data_nxt~0_combout ),
	.cout());
defparam \av_ld_aligning_data_nxt~0 .lut_mask = 16'hBEFF;
defparam \av_ld_aligning_data_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_aligning_data_nxt~1 (
	.dataa(d_read1),
	.datab(gnd),
	.datac(WideOr1),
	.datad(WideOr13),
	.cin(gnd),
	.combout(\av_ld_aligning_data_nxt~1_combout ),
	.cout());
defparam \av_ld_aligning_data_nxt~1 .lut_mask = 16'hAFFF;
defparam \av_ld_aligning_data_nxt~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_mem32~0 (
	.dataa(\D_iw[0]~q ),
	.datab(\D_iw[2]~q ),
	.datac(\D_iw[4]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\D_ctrl_mem32~0_combout ),
	.cout());
defparam \D_ctrl_mem32~0 .lut_mask = 16'hFEFF;
defparam \D_ctrl_mem32~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \av_ld_aligning_data_nxt~2 (
	.dataa(\av_ld_aligning_data_nxt~0_combout ),
	.datab(\av_ld_aligning_data_nxt~1_combout ),
	.datac(\av_ld_aligning_data~q ),
	.datad(\D_ctrl_mem32~0_combout ),
	.cin(gnd),
	.combout(\av_ld_aligning_data_nxt~2_combout ),
	.cout());
defparam \av_ld_aligning_data_nxt~2 .lut_mask = 16'hEFFF;
defparam \av_ld_aligning_data_nxt~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_stall~3 (
	.dataa(\E_valid_from_R~q ),
	.datab(\av_ld_waiting_for_data_nxt~1_combout ),
	.datac(\av_ld_aligning_data_nxt~2_combout ),
	.datad(\D_ctrl_mem32~0_combout ),
	.cin(gnd),
	.combout(\E_stall~3_combout ),
	.cout());
defparam \E_stall~3 .lut_mask = 16'hFEFF;
defparam \E_stall~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_stall~4 (
	.dataa(\E_new_inst~q ),
	.datab(\R_ctrl_st~q ),
	.datac(\R_ctrl_ld~q ),
	.datad(\E_stall~3_combout ),
	.cin(gnd),
	.combout(\E_stall~4_combout ),
	.cout());
defparam \E_stall~4 .lut_mask = 16'hFFFE;
defparam \E_stall~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_stall~5 (
	.dataa(d_write1),
	.datab(av_waitrequest),
	.datac(\E_stall~2_combout ),
	.datad(\E_stall~4_combout ),
	.cin(gnd),
	.combout(\E_stall~5_combout ),
	.cout());
defparam \E_stall~5 .lut_mask = 16'hFFFE;
defparam \E_stall~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_valid_from_R~0 (
	.dataa(\R_valid~q ),
	.datab(\E_stall~5_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\E_valid_from_R~0_combout ),
	.cout());
defparam \E_valid_from_R~0 .lut_mask = 16'hEEEE;
defparam \E_valid_from_R~0 .sum_lutc_input = "datac";

dffeas E_valid_from_R(
	.clk(clk_clk),
	.d(\E_valid_from_R~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_valid_from_R~q ),
	.prn(vcc));
defparam E_valid_from_R.is_wysiwyg = "true";
defparam E_valid_from_R.power_up = "low";

cycloneive_lcell_comb \W_valid~0 (
	.dataa(\E_valid_from_R~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\E_stall~5_combout ),
	.cin(gnd),
	.combout(\W_valid~0_combout ),
	.cout());
defparam \W_valid~0 .lut_mask = 16'hAAFF;
defparam \W_valid~0 .sum_lutc_input = "datac";

dffeas W_valid(
	.clk(clk_clk),
	.d(\W_valid~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_valid~q ),
	.prn(vcc));
defparam W_valid.is_wysiwyg = "true";
defparam W_valid.power_up = "low";

cycloneive_lcell_comb \hbreak_pending_nxt~0 (
	.dataa(\hbreak_pending~q ),
	.datab(\hbreak_req~0_combout ),
	.datac(gnd),
	.datad(hbreak_enabled1),
	.cin(gnd),
	.combout(\hbreak_pending_nxt~0_combout ),
	.cout());
defparam \hbreak_pending_nxt~0 .lut_mask = 16'hEEFF;
defparam \hbreak_pending_nxt~0 .sum_lutc_input = "datac";

dffeas hbreak_pending(
	.clk(clk_clk),
	.d(\hbreak_pending_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\hbreak_pending~q ),
	.prn(vcc));
defparam hbreak_pending.is_wysiwyg = "true";
defparam hbreak_pending.power_up = "low";

cycloneive_lcell_comb \wait_for_one_post_bret_inst~0 (
	.dataa(\the_nios_mcu_nios_cpu_cpu_nios2_oci|the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_single_step_mode~q ),
	.datab(hbreak_enabled1),
	.datac(\wait_for_one_post_bret_inst~q ),
	.datad(\F_valid~0_combout ),
	.cin(gnd),
	.combout(\wait_for_one_post_bret_inst~0_combout ),
	.cout());
defparam \wait_for_one_post_bret_inst~0 .lut_mask = 16'hFEFF;
defparam \wait_for_one_post_bret_inst~0 .sum_lutc_input = "datac";

dffeas wait_for_one_post_bret_inst(
	.clk(clk_clk),
	.d(\wait_for_one_post_bret_inst~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wait_for_one_post_bret_inst~q ),
	.prn(vcc));
defparam wait_for_one_post_bret_inst.is_wysiwyg = "true";
defparam wait_for_one_post_bret_inst.power_up = "low";

cycloneive_lcell_comb \hbreak_req~0 (
	.dataa(\W_valid~q ),
	.datab(\hbreak_pending~q ),
	.datac(\the_nios_mcu_nios_cpu_cpu_nios2_oci|the_nios_mcu_nios_cpu_cpu_nios2_oci_debug|jtag_break~q ),
	.datad(\wait_for_one_post_bret_inst~q ),
	.cin(gnd),
	.combout(\hbreak_req~0_combout ),
	.cout());
defparam \hbreak_req~0 .lut_mask = 16'hFEFF;
defparam \hbreak_req~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_jmp_direct~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\D_iw[5]~q ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_jmp_direct~0_combout ),
	.cout());
defparam \D_ctrl_jmp_direct~0 .lut_mask = 16'h0FFF;
defparam \D_ctrl_jmp_direct~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_jmp_direct~1 (
	.dataa(\D_ctrl_jmp_direct~0_combout ),
	.datab(\D_iw[1]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\D_ctrl_jmp_direct~1_combout ),
	.cout());
defparam \D_ctrl_jmp_direct~1 .lut_mask = 16'hBFFF;
defparam \D_ctrl_jmp_direct~1 .sum_lutc_input = "datac";

dffeas R_ctrl_jmp_direct(
	.clk(clk_clk),
	.d(\D_ctrl_jmp_direct~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_jmp_direct~q ),
	.prn(vcc));
defparam R_ctrl_jmp_direct.is_wysiwyg = "true";
defparam R_ctrl_jmp_direct.power_up = "low";

dffeas R_ctrl_br(
	.clk(clk_clk),
	.d(\R_ctrl_br_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_br~q ),
	.prn(vcc));
defparam R_ctrl_br.is_wysiwyg = "true";
defparam R_ctrl_br.power_up = "low";

cycloneive_lcell_comb \D_ctrl_retaddr~3 (
	.dataa(\Equal62~13_combout ),
	.datab(\Equal62~12_combout ),
	.datac(\D_iw[15]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~3_combout ),
	.cout());
defparam \D_ctrl_retaddr~3 .lut_mask = 16'hEFFF;
defparam \D_ctrl_retaddr~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_retaddr~4 (
	.dataa(\D_ctrl_retaddr~3_combout ),
	.datab(\Equal62~8_combout ),
	.datac(\Equal62~14_combout ),
	.datad(\D_ctrl_implicit_dst_eretaddr~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~4_combout ),
	.cout());
defparam \D_ctrl_retaddr~4 .lut_mask = 16'hFEFF;
defparam \D_ctrl_retaddr~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_retaddr~5 (
	.dataa(\Equal0~7_combout ),
	.datab(\D_ctrl_retaddr~4_combout ),
	.datac(\D_ctrl_force_src2_zero~6_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~5_combout ),
	.cout());
defparam \D_ctrl_retaddr~5 .lut_mask = 16'hF7F7;
defparam \D_ctrl_retaddr~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~9 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~9_combout ),
	.cout());
defparam \Equal0~9 .lut_mask = 16'hFF7F;
defparam \Equal0~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_retaddr~6 (
	.dataa(\Equal0~12_combout ),
	.datab(\D_ctrl_force_src2_zero~0_combout ),
	.datac(\Equal0~9_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~6_combout ),
	.cout());
defparam \D_ctrl_retaddr~6 .lut_mask = 16'hFDFE;
defparam \D_ctrl_retaddr~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_retaddr~7 (
	.dataa(\D_iw[5]~q ),
	.datab(\Equal0~16_combout ),
	.datac(\D_iw[4]~q ),
	.datad(\D_ctrl_retaddr~6_combout ),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~7_combout ),
	.cout());
defparam \D_ctrl_retaddr~7 .lut_mask = 16'hFFBE;
defparam \D_ctrl_retaddr~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_retaddr~8 (
	.dataa(\Equal0~2_combout ),
	.datab(\D_ctrl_retaddr~5_combout ),
	.datac(\D_iw[4]~q ),
	.datad(\D_ctrl_retaddr~7_combout ),
	.cin(gnd),
	.combout(\D_ctrl_retaddr~8_combout ),
	.cout());
defparam \D_ctrl_retaddr~8 .lut_mask = 16'hBFFB;
defparam \D_ctrl_retaddr~8 .sum_lutc_input = "datac";

dffeas R_ctrl_retaddr(
	.clk(clk_clk),
	.d(\D_ctrl_retaddr~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_retaddr~q ),
	.prn(vcc));
defparam R_ctrl_retaddr.is_wysiwyg = "true";
defparam R_ctrl_retaddr.power_up = "low";

cycloneive_lcell_comb \R_src1~37 (
	.dataa(\R_valid~q ),
	.datab(\E_valid_from_R~q ),
	.datac(\R_ctrl_br~q ),
	.datad(\R_ctrl_retaddr~q ),
	.cin(gnd),
	.combout(\R_src1~37_combout ),
	.cout());
defparam \R_src1~37 .lut_mask = 16'hFFFE;
defparam \R_src1~37 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src1[0]~39 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[0] ),
	.datad(\R_src1~37_combout ),
	.cin(gnd),
	.combout(\R_src1[0]~39_combout ),
	.cout());
defparam \R_src1[0]~39 .lut_mask = 16'hF7FF;
defparam \R_src1[0]~39 .sum_lutc_input = "datac";

dffeas \E_src1[0] (
	.clk(clk_clk),
	.d(\R_src1[0]~39_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[0]~q ),
	.prn(vcc));
defparam \E_src1[0] .is_wysiwyg = "true";
defparam \E_src1[0] .power_up = "low";

cycloneive_lcell_comb D_op_wrctl(
	.dataa(\Equal0~7_combout ),
	.datab(\D_iw[14]~q ),
	.datac(\Equal62~3_combout ),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_op_wrctl~combout ),
	.cout());
defparam D_op_wrctl.lut_mask = 16'hFEFF;
defparam D_op_wrctl.sum_lutc_input = "datac";

dffeas R_ctrl_wrctl_inst(
	.clk(clk_clk),
	.d(\D_op_wrctl~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_wrctl_inst~q ),
	.prn(vcc));
defparam R_ctrl_wrctl_inst.is_wysiwyg = "true";
defparam R_ctrl_wrctl_inst.power_up = "low";

cycloneive_lcell_comb \E_wrctl_status~0 (
	.dataa(\R_ctrl_wrctl_inst~q ),
	.datab(\D_iw[10]~q ),
	.datac(\D_iw[8]~q ),
	.datad(\D_iw[9]~q ),
	.cin(gnd),
	.combout(\E_wrctl_status~0_combout ),
	.cout());
defparam \E_wrctl_status~0 .lut_mask = 16'hBFFF;
defparam \E_wrctl_status~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_estatus_reg_inst_nxt~0 (
	.dataa(\E_src1[0]~q ),
	.datab(\D_iw[6]~q ),
	.datac(\E_wrctl_status~0_combout ),
	.datad(\D_iw[7]~q ),
	.cin(gnd),
	.combout(\W_estatus_reg_inst_nxt~0_combout ),
	.cout());
defparam \W_estatus_reg_inst_nxt~0 .lut_mask = 16'hFEFF;
defparam \W_estatus_reg_inst_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_estatus_reg_inst_nxt~1 (
	.dataa(\W_estatus_reg~q ),
	.datab(\D_iw[7]~q ),
	.datac(\D_iw[6]~q ),
	.datad(\E_wrctl_status~0_combout ),
	.cin(gnd),
	.combout(\W_estatus_reg_inst_nxt~1_combout ),
	.cout());
defparam \W_estatus_reg_inst_nxt~1 .lut_mask = 16'hEFFF;
defparam \W_estatus_reg_inst_nxt~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~3 (
	.dataa(\D_op_opx_rsv63~0_combout ),
	.datab(\Equal62~14_combout ),
	.datac(\Equal62~8_combout ),
	.datad(\D_ctrl_implicit_dst_eretaddr~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~3_combout ),
	.cout());
defparam \D_ctrl_exception~3 .lut_mask = 16'hFEFF;
defparam \D_ctrl_exception~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_implicit_dst_eretaddr~16 (
	.dataa(\D_iw[16]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~16_combout ),
	.cout());
defparam \D_ctrl_implicit_dst_eretaddr~16 .lut_mask = 16'hAAFF;
defparam \D_ctrl_implicit_dst_eretaddr~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~4 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[12]~q ),
	.datac(\D_iw[13]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_ctrl_exception~4_combout ),
	.cout());
defparam \D_ctrl_exception~4 .lut_mask = 16'hFBFF;
defparam \D_ctrl_exception~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~5 (
	.dataa(\Equal0~7_combout ),
	.datab(\D_ctrl_exception~3_combout ),
	.datac(\D_ctrl_implicit_dst_eretaddr~16_combout ),
	.datad(\D_ctrl_exception~4_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~5_combout ),
	.cout());
defparam \D_ctrl_exception~5 .lut_mask = 16'hFFFE;
defparam \D_ctrl_exception~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_implicit_dst_eretaddr~13 (
	.dataa(\D_ctrl_implicit_dst_eretaddr~5_combout ),
	.datab(\D_ctrl_implicit_dst_eretaddr~10_combout ),
	.datac(\D_ctrl_implicit_dst_eretaddr~12_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~13_combout ),
	.cout());
defparam \D_ctrl_implicit_dst_eretaddr~13 .lut_mask = 16'hFEFE;
defparam \D_ctrl_implicit_dst_eretaddr~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~0 (
	.dataa(\D_iw[5]~q ),
	.datab(\Equal0~12_combout ),
	.datac(\Equal0~9_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_exception~0_combout ),
	.cout());
defparam \D_ctrl_exception~0 .lut_mask = 16'hFEFF;
defparam \D_ctrl_exception~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~1 (
	.dataa(\Equal0~3_combout ),
	.datab(\Equal0~2_combout ),
	.datac(\Equal0~16_combout ),
	.datad(\D_ctrl_exception~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~1_combout ),
	.cout());
defparam \D_ctrl_exception~1 .lut_mask = 16'hBFFF;
defparam \D_ctrl_exception~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~2 (
	.dataa(\D_ctrl_exception~1_combout ),
	.datab(\D_ctrl_force_src2_zero~0_combout ),
	.datac(\Equal0~12_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_exception~2_combout ),
	.cout());
defparam \D_ctrl_exception~2 .lut_mask = 16'hEFFF;
defparam \D_ctrl_exception~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_exception~6 (
	.dataa(\D_ctrl_exception~5_combout ),
	.datab(gnd),
	.datac(\D_ctrl_implicit_dst_eretaddr~13_combout ),
	.datad(\D_ctrl_exception~2_combout ),
	.cin(gnd),
	.combout(\D_ctrl_exception~6_combout ),
	.cout());
defparam \D_ctrl_exception~6 .lut_mask = 16'hAFFF;
defparam \D_ctrl_exception~6 .sum_lutc_input = "datac";

dffeas R_ctrl_exception(
	.clk(clk_clk),
	.d(\D_ctrl_exception~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_exception~q ),
	.prn(vcc));
defparam R_ctrl_exception.is_wysiwyg = "true";
defparam R_ctrl_exception.power_up = "low";

cycloneive_lcell_comb \W_estatus_reg_inst_nxt~2 (
	.dataa(\W_status_reg_pie~q ),
	.datab(\W_estatus_reg_inst_nxt~0_combout ),
	.datac(\W_estatus_reg_inst_nxt~1_combout ),
	.datad(\R_ctrl_exception~q ),
	.cin(gnd),
	.combout(\W_estatus_reg_inst_nxt~2_combout ),
	.cout());
defparam \W_estatus_reg_inst_nxt~2 .lut_mask = 16'hFAFC;
defparam \W_estatus_reg_inst_nxt~2 .sum_lutc_input = "datac";

dffeas W_estatus_reg(
	.clk(clk_clk),
	.d(\W_estatus_reg_inst_nxt~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\E_valid_from_R~q ),
	.q(\W_estatus_reg~q ),
	.prn(vcc));
defparam W_estatus_reg.is_wysiwyg = "true";
defparam W_estatus_reg.power_up = "low";

cycloneive_lcell_comb \W_bstatus_reg_inst_nxt~0 (
	.dataa(\E_src1[0]~q ),
	.datab(\D_iw[7]~q ),
	.datac(\E_wrctl_status~0_combout ),
	.datad(\D_iw[6]~q ),
	.cin(gnd),
	.combout(\W_bstatus_reg_inst_nxt~0_combout ),
	.cout());
defparam \W_bstatus_reg_inst_nxt~0 .lut_mask = 16'hFEFF;
defparam \W_bstatus_reg_inst_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_bstatus_reg_inst_nxt~1 (
	.dataa(\W_bstatus_reg~q ),
	.datab(\D_iw[6]~q ),
	.datac(\D_iw[7]~q ),
	.datad(\E_wrctl_status~0_combout ),
	.cin(gnd),
	.combout(\W_bstatus_reg_inst_nxt~1_combout ),
	.cout());
defparam \W_bstatus_reg_inst_nxt~1 .lut_mask = 16'hEFFF;
defparam \W_bstatus_reg_inst_nxt~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_break~0 (
	.dataa(\D_iw[13]~q ),
	.datab(\D_iw[16]~q ),
	.datac(\D_op_opx_rsv17~0_combout ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\D_ctrl_break~0_combout ),
	.cout());
defparam \D_ctrl_break~0 .lut_mask = 16'hFEFF;
defparam \D_ctrl_break~0 .sum_lutc_input = "datac";

dffeas R_ctrl_break(
	.clk(clk_clk),
	.d(\D_ctrl_break~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_break~q ),
	.prn(vcc));
defparam R_ctrl_break.is_wysiwyg = "true";
defparam R_ctrl_break.power_up = "low";

cycloneive_lcell_comb \W_bstatus_reg_inst_nxt~2 (
	.dataa(\W_status_reg_pie~q ),
	.datab(\W_bstatus_reg_inst_nxt~0_combout ),
	.datac(\W_bstatus_reg_inst_nxt~1_combout ),
	.datad(\R_ctrl_break~q ),
	.cin(gnd),
	.combout(\W_bstatus_reg_inst_nxt~2_combout ),
	.cout());
defparam \W_bstatus_reg_inst_nxt~2 .lut_mask = 16'hFAFC;
defparam \W_bstatus_reg_inst_nxt~2 .sum_lutc_input = "datac";

dffeas W_bstatus_reg(
	.clk(clk_clk),
	.d(\W_bstatus_reg_inst_nxt~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\E_valid_from_R~q ),
	.q(\W_bstatus_reg~q ),
	.prn(vcc));
defparam W_bstatus_reg.is_wysiwyg = "true";
defparam W_bstatus_reg.power_up = "low";

cycloneive_lcell_comb \E_wrctl_status~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\D_iw[7]~q ),
	.datad(\D_iw[6]~q ),
	.cin(gnd),
	.combout(\E_wrctl_status~1_combout ),
	.cout());
defparam \E_wrctl_status~1 .lut_mask = 16'h0FFF;
defparam \E_wrctl_status~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_status_reg_pie_inst_nxt~0 (
	.dataa(\E_src1[0]~q ),
	.datab(\W_status_reg_pie~q ),
	.datac(\E_wrctl_status~1_combout ),
	.datad(\E_wrctl_status~0_combout ),
	.cin(gnd),
	.combout(\W_status_reg_pie_inst_nxt~0_combout ),
	.cout());
defparam \W_status_reg_pie_inst_nxt~0 .lut_mask = 16'hEFFE;
defparam \W_status_reg_pie_inst_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_status_reg_pie_inst_nxt~1 (
	.dataa(\W_bstatus_reg~q ),
	.datab(\W_status_reg_pie_inst_nxt~0_combout ),
	.datac(\D_op_cmpge~0_combout ),
	.datad(\Equal62~9_combout ),
	.cin(gnd),
	.combout(\W_status_reg_pie_inst_nxt~1_combout ),
	.cout());
defparam \W_status_reg_pie_inst_nxt~1 .lut_mask = 16'hEFFE;
defparam \W_status_reg_pie_inst_nxt~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb D_op_eret(
	.dataa(\Equal0~7_combout ),
	.datab(\Equal62~9_combout ),
	.datac(\D_iw[15]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_op_eret~combout ),
	.cout());
defparam D_op_eret.lut_mask = 16'hEFFF;
defparam D_op_eret.sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_sel_nxt.10~0 (
	.dataa(\R_ctrl_exception~q ),
	.datab(\R_ctrl_break~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\F_pc_sel_nxt.10~0_combout ),
	.cout());
defparam \F_pc_sel_nxt.10~0 .lut_mask = 16'hEEEE;
defparam \F_pc_sel_nxt.10~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_status_reg_pie_inst_nxt~2 (
	.dataa(\W_estatus_reg~q ),
	.datab(\W_status_reg_pie_inst_nxt~1_combout ),
	.datac(\D_op_eret~combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\W_status_reg_pie_inst_nxt~2_combout ),
	.cout());
defparam \W_status_reg_pie_inst_nxt~2 .lut_mask = 16'hACFF;
defparam \W_status_reg_pie_inst_nxt~2 .sum_lutc_input = "datac";

dffeas W_status_reg_pie(
	.clk(clk_clk),
	.d(\W_status_reg_pie_inst_nxt~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\E_valid_from_R~q ),
	.q(\W_status_reg_pie~q ),
	.prn(vcc));
defparam W_status_reg_pie.is_wysiwyg = "true";
defparam W_status_reg_pie.power_up = "low";

cycloneive_lcell_comb \W_ienable_reg_nxt~0 (
	.dataa(\E_valid_from_R~q ),
	.datab(\D_iw[7]~q ),
	.datac(\D_iw[6]~q ),
	.datad(\E_wrctl_status~0_combout ),
	.cin(gnd),
	.combout(\W_ienable_reg_nxt~0_combout ),
	.cout());
defparam \W_ienable_reg_nxt~0 .lut_mask = 16'hFFFE;
defparam \W_ienable_reg_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_ienable_reg[0]~0 (
	.dataa(\E_src1[0]~q ),
	.datab(\W_ienable_reg[0]~q ),
	.datac(gnd),
	.datad(\W_ienable_reg_nxt~0_combout ),
	.cin(gnd),
	.combout(\W_ienable_reg[0]~0_combout ),
	.cout());
defparam \W_ienable_reg[0]~0 .lut_mask = 16'hAACC;
defparam \W_ienable_reg[0]~0 .sum_lutc_input = "datac";

dffeas \W_ienable_reg[0] (
	.clk(clk_clk),
	.d(\W_ienable_reg[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_ienable_reg[0]~q ),
	.prn(vcc));
defparam \W_ienable_reg[0] .is_wysiwyg = "true";
defparam \W_ienable_reg[0] .power_up = "low";

cycloneive_lcell_comb \W_ipending_reg_nxt[0]~0 (
	.dataa(\W_ienable_reg[0]~q ),
	.datab(av_readdata_9),
	.datac(av_readdata_8),
	.datad(\the_nios_mcu_nios_cpu_cpu_nios2_oci|the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_ienable[0]~q ),
	.cin(gnd),
	.combout(\W_ipending_reg_nxt[0]~0_combout ),
	.cout());
defparam \W_ipending_reg_nxt[0]~0 .lut_mask = 16'hFEFF;
defparam \W_ipending_reg_nxt[0]~0 .sum_lutc_input = "datac";

dffeas \W_ipending_reg[0] (
	.clk(clk_clk),
	.d(\W_ipending_reg_nxt[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_ipending_reg[0]~q ),
	.prn(vcc));
defparam \W_ipending_reg[0] .is_wysiwyg = "true";
defparam \W_ipending_reg[0] .power_up = "low";

cycloneive_lcell_comb \D_iw[27]~0 (
	.dataa(hbreak_enabled1),
	.datab(\hbreak_req~0_combout ),
	.datac(\W_status_reg_pie~q ),
	.datad(\W_ipending_reg[0]~q ),
	.cin(gnd),
	.combout(\D_iw[27]~0_combout ),
	.cout());
defparam \D_iw[27]~0 .lut_mask = 16'hBFFF;
defparam \D_iw[27]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[11]~10 (
	.dataa(src_payload),
	.datab(src1_valid),
	.datac(av_readdata_pre_11),
	.datad(\D_iw[27]~0_combout ),
	.cin(gnd),
	.combout(\F_iw[11]~10_combout ),
	.cout());
defparam \F_iw[11]~10 .lut_mask = 16'hFEFF;
defparam \F_iw[11]~10 .sum_lutc_input = "datac";

dffeas \D_iw[11] (
	.clk(clk_clk),
	.d(\F_iw[11]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[11]~q ),
	.prn(vcc));
defparam \D_iw[11] .is_wysiwyg = "true";
defparam \D_iw[11] .power_up = "low";

cycloneive_lcell_comb \Equal62~0 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[13]~q ),
	.datac(\D_iw[16]~q ),
	.datad(\D_iw[12]~q ),
	.cin(gnd),
	.combout(\Equal62~0_combout ),
	.cout());
defparam \Equal62~0 .lut_mask = 16'h7FFF;
defparam \Equal62~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~5 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~5_combout ),
	.cout());
defparam \Equal0~5 .lut_mask = 16'hFFBF;
defparam \Equal0~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_invert_arith_src_msb~0 (
	.dataa(\D_iw[4]~q ),
	.datab(\Equal0~4_combout ),
	.datac(\Equal0~5_combout ),
	.datad(\D_ctrl_alu_force_xor~14_combout ),
	.cin(gnd),
	.combout(\E_invert_arith_src_msb~0_combout ),
	.cout());
defparam \E_invert_arith_src_msb~0 .lut_mask = 16'h27FF;
defparam \E_invert_arith_src_msb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_alu_subtract~2 (
	.dataa(\Equal62~0_combout ),
	.datab(\D_op_cmpge~0_combout ),
	.datac(gnd),
	.datad(\E_invert_arith_src_msb~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_alu_subtract~2_combout ),
	.cout());
defparam \D_ctrl_alu_subtract~2 .lut_mask = 16'hEEFF;
defparam \D_ctrl_alu_subtract~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_alu_subtract~3 (
	.dataa(\Equal62~2_combout ),
	.datab(\Equal62~1_combout ),
	.datac(\Equal62~0_combout ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_ctrl_alu_subtract~3_combout ),
	.cout());
defparam \D_ctrl_alu_subtract~3 .lut_mask = 16'hFAFC;
defparam \D_ctrl_alu_subtract~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_alu_subtract~4 (
	.dataa(\D_iw[14]~q ),
	.datab(\D_iw[15]~q ),
	.datac(\Equal62~1_combout ),
	.datad(\D_ctrl_alu_subtract~3_combout ),
	.cin(gnd),
	.combout(\D_ctrl_alu_subtract~4_combout ),
	.cout());
defparam \D_ctrl_alu_subtract~4 .lut_mask = 16'hFFB8;
defparam \D_ctrl_alu_subtract~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_alu_sub~0 (
	.dataa(\R_valid~q ),
	.datab(\D_ctrl_alu_subtract~2_combout ),
	.datac(\Equal0~7_combout ),
	.datad(\D_ctrl_alu_subtract~4_combout ),
	.cin(gnd),
	.combout(\E_alu_sub~0_combout ),
	.cout());
defparam \E_alu_sub~0 .lut_mask = 16'hFFFE;
defparam \E_alu_sub~0 .sum_lutc_input = "datac";

dffeas E_alu_sub(
	.clk(clk_clk),
	.d(\E_alu_sub~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_alu_sub~q ),
	.prn(vcc));
defparam E_alu_sub.is_wysiwyg = "true";
defparam E_alu_sub.power_up = "low";

cycloneive_lcell_comb \F_iw[18]~26 (
	.dataa(src1_valid),
	.datab(read_latency_shift_reg_05),
	.datac(q_a_18),
	.datad(av_readdata_pre_18),
	.cin(gnd),
	.combout(\F_iw[18]~26_combout ),
	.cout());
defparam \F_iw[18]~26 .lut_mask = 16'hFFFE;
defparam \F_iw[18]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[18]~27 (
	.dataa(\D_iw[27]~0_combout ),
	.datab(\F_iw[18]~26_combout ),
	.datac(\hbreak_req~0_combout ),
	.datad(hbreak_enabled1),
	.cin(gnd),
	.combout(\F_iw[18]~27_combout ),
	.cout());
defparam \F_iw[18]~27 .lut_mask = 16'hFEFF;
defparam \F_iw[18]~27 .sum_lutc_input = "datac";

dffeas \D_iw[18] (
	.clk(clk_clk),
	.d(\F_iw[18]~27_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[18]~q ),
	.prn(vcc));
defparam \D_iw[18] .is_wysiwyg = "true";
defparam \D_iw[18] .power_up = "low";

cycloneive_lcell_comb \E_src2[7]~15 (
	.dataa(\R_ctrl_src_imm5_shift_rot~q ),
	.datab(\R_ctrl_hi_imm16~q ),
	.datac(\R_ctrl_force_src2_zero~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\E_src2[7]~15_combout ),
	.cout());
defparam \E_src2[7]~15 .lut_mask = 16'hFEFE;
defparam \E_src2[7]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_lo[12]~0 (
	.dataa(\D_iw[18]~q ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[7]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[12]~0_combout ),
	.cout());
defparam \R_src2_lo[12]~0 .lut_mask = 16'hACFF;
defparam \R_src2_lo[12]~0 .sum_lutc_input = "datac";

dffeas \E_src2[12] (
	.clk(clk_clk),
	.d(\R_src2_lo[12]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[12]~q ),
	.prn(vcc));
defparam \E_src2[12] .is_wysiwyg = "true";
defparam \E_src2[12] .power_up = "low";

cycloneive_lcell_comb \Add1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[12]~q ),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout());
defparam \Add1~0 .lut_mask = 16'h0FF0;
defparam \Add1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src1~36 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_valid_from_R~q ),
	.datad(\R_ctrl_jmp_direct~q ),
	.cin(gnd),
	.combout(\R_src1~36_combout ),
	.cout());
defparam \R_src1~36 .lut_mask = 16'h0FFF;
defparam \R_src1~36 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[12]~3 (
	.dataa(\D_iw[16]~q ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[12] ),
	.datac(gnd),
	.datad(\R_src1~36_combout ),
	.cin(gnd),
	.combout(\E_src1[12]~3_combout ),
	.cout());
defparam \E_src1[12]~3 .lut_mask = 16'hAACC;
defparam \E_src1[12]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_plus_one[0]~0 (
	.dataa(F_pc_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\F_pc_plus_one[0]~0_combout ),
	.cout(\F_pc_plus_one[0]~1 ));
defparam \F_pc_plus_one[0]~0 .lut_mask = 16'h55AA;
defparam \F_pc_plus_one[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_plus_one[1]~2 (
	.dataa(F_pc_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[0]~1 ),
	.combout(\F_pc_plus_one[1]~2_combout ),
	.cout(\F_pc_plus_one[1]~3 ));
defparam \F_pc_plus_one[1]~2 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[1]~2 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[2]~4 (
	.dataa(F_pc_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[1]~3 ),
	.combout(\F_pc_plus_one[2]~4_combout ),
	.cout(\F_pc_plus_one[2]~5 ));
defparam \F_pc_plus_one[2]~4 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[2]~4 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[3]~6 (
	.dataa(F_pc_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[2]~5 ),
	.combout(\F_pc_plus_one[3]~6_combout ),
	.cout(\F_pc_plus_one[3]~7 ));
defparam \F_pc_plus_one[3]~6 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[3]~6 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[4]~8 (
	.dataa(F_pc_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[3]~7 ),
	.combout(\F_pc_plus_one[4]~8_combout ),
	.cout(\F_pc_plus_one[4]~9 ));
defparam \F_pc_plus_one[4]~8 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[4]~8 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[5]~10 (
	.dataa(F_pc_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[4]~9 ),
	.combout(\F_pc_plus_one[5]~10_combout ),
	.cout(\F_pc_plus_one[5]~11 ));
defparam \F_pc_plus_one[5]~10 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[5]~10 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[6]~12 (
	.dataa(F_pc_6),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[5]~11 ),
	.combout(\F_pc_plus_one[6]~12_combout ),
	.cout(\F_pc_plus_one[6]~13 ));
defparam \F_pc_plus_one[6]~12 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[6]~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[7]~14 (
	.dataa(F_pc_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[6]~13 ),
	.combout(\F_pc_plus_one[7]~14_combout ),
	.cout(\F_pc_plus_one[7]~15 ));
defparam \F_pc_plus_one[7]~14 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[7]~14 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[8]~16 (
	.dataa(F_pc_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[7]~15 ),
	.combout(\F_pc_plus_one[8]~16_combout ),
	.cout(\F_pc_plus_one[8]~17 ));
defparam \F_pc_plus_one[8]~16 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[8]~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[9]~18 (
	.dataa(F_pc_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[8]~17 ),
	.combout(\F_pc_plus_one[9]~18_combout ),
	.cout(\F_pc_plus_one[9]~19 ));
defparam \F_pc_plus_one[9]~18 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[9]~18 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[10]~20 (
	.dataa(F_pc_10),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[9]~19 ),
	.combout(\F_pc_plus_one[10]~20_combout ),
	.cout(\F_pc_plus_one[10]~21 ));
defparam \F_pc_plus_one[10]~20 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[10]~20 .sum_lutc_input = "cin";

dffeas \E_src1[12] (
	.clk(clk_clk),
	.d(\E_src1[12]~3_combout ),
	.asdata(\F_pc_plus_one[10]~20_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~37_combout ),
	.ena(vcc),
	.q(\E_src1[12]~q ),
	.prn(vcc));
defparam \E_src1[12] .is_wysiwyg = "true";
defparam \E_src1[12] .power_up = "low";

cycloneive_lcell_comb \F_iw[17]~28 (
	.dataa(src1_valid),
	.datab(read_latency_shift_reg_05),
	.datac(q_a_17),
	.datad(av_readdata_pre_17),
	.cin(gnd),
	.combout(\F_iw[17]~28_combout ),
	.cout());
defparam \F_iw[17]~28 .lut_mask = 16'hFFFE;
defparam \F_iw[17]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[17]~29 (
	.dataa(\F_iw[17]~28_combout ),
	.datab(hbreak_enabled1),
	.datac(\hbreak_req~0_combout ),
	.datad(\D_iw[27]~0_combout ),
	.cin(gnd),
	.combout(\F_iw[17]~29_combout ),
	.cout());
defparam \F_iw[17]~29 .lut_mask = 16'hAFCF;
defparam \F_iw[17]~29 .sum_lutc_input = "datac";

dffeas \D_iw[17] (
	.clk(clk_clk),
	.d(\F_iw[17]~29_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[17]~q ),
	.prn(vcc));
defparam \D_iw[17] .is_wysiwyg = "true";
defparam \D_iw[17] .power_up = "low";

cycloneive_lcell_comb \R_src2_lo[11]~1 (
	.dataa(\D_iw[17]~q ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[7]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[11]~1_combout ),
	.cout());
defparam \R_src2_lo[11]~1 .lut_mask = 16'hACFF;
defparam \R_src2_lo[11]~1 .sum_lutc_input = "datac";

dffeas \E_src2[11] (
	.clk(clk_clk),
	.d(\R_src2_lo[11]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[11]~q ),
	.prn(vcc));
defparam \E_src2[11] .is_wysiwyg = "true";
defparam \E_src2[11] .power_up = "low";

cycloneive_lcell_comb \Add1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[11]~q ),
	.cin(gnd),
	.combout(\Add1~1_combout ),
	.cout());
defparam \Add1~1 .lut_mask = 16'h0FF0;
defparam \Add1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[11]~4 (
	.dataa(\D_iw[15]~q ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[11] ),
	.datac(gnd),
	.datad(\R_src1~36_combout ),
	.cin(gnd),
	.combout(\E_src1[11]~4_combout ),
	.cout());
defparam \E_src1[11]~4 .lut_mask = 16'hAACC;
defparam \E_src1[11]~4 .sum_lutc_input = "datac";

dffeas \E_src1[11] (
	.clk(clk_clk),
	.d(\E_src1[11]~4_combout ),
	.asdata(\F_pc_plus_one[9]~18_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~37_combout ),
	.ena(vcc),
	.q(\E_src1[11]~q ),
	.prn(vcc));
defparam \E_src1[11] .is_wysiwyg = "true";
defparam \E_src1[11] .power_up = "low";

cycloneive_lcell_comb \R_src2_lo[10]~2 (
	.dataa(\D_iw[16]~q ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[7]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[10]~2_combout ),
	.cout());
defparam \R_src2_lo[10]~2 .lut_mask = 16'hACFF;
defparam \R_src2_lo[10]~2 .sum_lutc_input = "datac";

dffeas \E_src2[10] (
	.clk(clk_clk),
	.d(\R_src2_lo[10]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[10]~q ),
	.prn(vcc));
defparam \E_src2[10] .is_wysiwyg = "true";
defparam \E_src2[10] .power_up = "low";

cycloneive_lcell_comb \Add1~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[10]~q ),
	.cin(gnd),
	.combout(\Add1~2_combout ),
	.cout());
defparam \Add1~2 .lut_mask = 16'h0FF0;
defparam \Add1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[10]~5 (
	.dataa(\D_iw[14]~q ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[10] ),
	.datac(gnd),
	.datad(\R_src1~36_combout ),
	.cin(gnd),
	.combout(\E_src1[10]~5_combout ),
	.cout());
defparam \E_src1[10]~5 .lut_mask = 16'hAACC;
defparam \E_src1[10]~5 .sum_lutc_input = "datac";

dffeas \E_src1[10] (
	.clk(clk_clk),
	.d(\E_src1[10]~5_combout ),
	.asdata(\F_pc_plus_one[8]~16_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~37_combout ),
	.ena(vcc),
	.q(\E_src1[10]~q ),
	.prn(vcc));
defparam \E_src1[10] .is_wysiwyg = "true";
defparam \E_src1[10] .power_up = "low";

cycloneive_lcell_comb \R_src2_lo[9]~3 (
	.dataa(\D_iw[15]~q ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[7]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[9]~3_combout ),
	.cout());
defparam \R_src2_lo[9]~3 .lut_mask = 16'hACFF;
defparam \R_src2_lo[9]~3 .sum_lutc_input = "datac";

dffeas \E_src2[9] (
	.clk(clk_clk),
	.d(\R_src2_lo[9]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[9]~q ),
	.prn(vcc));
defparam \E_src2[9] .is_wysiwyg = "true";
defparam \E_src2[9] .power_up = "low";

cycloneive_lcell_comb \Add1~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[9]~q ),
	.cin(gnd),
	.combout(\Add1~3_combout ),
	.cout());
defparam \Add1~3 .lut_mask = 16'h0FF0;
defparam \Add1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[9]~6 (
	.dataa(\D_iw[13]~q ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[9] ),
	.datac(gnd),
	.datad(\R_src1~36_combout ),
	.cin(gnd),
	.combout(\E_src1[9]~6_combout ),
	.cout());
defparam \E_src1[9]~6 .lut_mask = 16'hAACC;
defparam \E_src1[9]~6 .sum_lutc_input = "datac";

dffeas \E_src1[9] (
	.clk(clk_clk),
	.d(\E_src1[9]~6_combout ),
	.asdata(\F_pc_plus_one[7]~14_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~37_combout ),
	.ena(vcc),
	.q(\E_src1[9]~q ),
	.prn(vcc));
defparam \E_src1[9] .is_wysiwyg = "true";
defparam \E_src1[9] .power_up = "low";

cycloneive_lcell_comb \R_src2_lo[8]~4 (
	.dataa(\D_iw[14]~q ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[7]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[8]~4_combout ),
	.cout());
defparam \R_src2_lo[8]~4 .lut_mask = 16'hACFF;
defparam \R_src2_lo[8]~4 .sum_lutc_input = "datac";

dffeas \E_src2[8] (
	.clk(clk_clk),
	.d(\R_src2_lo[8]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[8]~q ),
	.prn(vcc));
defparam \E_src2[8] .is_wysiwyg = "true";
defparam \E_src2[8] .power_up = "low";

cycloneive_lcell_comb \Add1~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[8]~q ),
	.cin(gnd),
	.combout(\Add1~4_combout ),
	.cout());
defparam \Add1~4 .lut_mask = 16'h0FF0;
defparam \Add1~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[8]~7 (
	.dataa(\D_iw[12]~q ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[8] ),
	.datac(gnd),
	.datad(\R_src1~36_combout ),
	.cin(gnd),
	.combout(\E_src1[8]~7_combout ),
	.cout());
defparam \E_src1[8]~7 .lut_mask = 16'hAACC;
defparam \E_src1[8]~7 .sum_lutc_input = "datac";

dffeas \E_src1[8] (
	.clk(clk_clk),
	.d(\E_src1[8]~7_combout ),
	.asdata(\F_pc_plus_one[6]~12_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~37_combout ),
	.ena(vcc),
	.q(\E_src1[8]~q ),
	.prn(vcc));
defparam \E_src1[8] .is_wysiwyg = "true";
defparam \E_src1[8] .power_up = "low";

cycloneive_lcell_comb \R_src2_lo[7]~5 (
	.dataa(\D_iw[13]~q ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[7]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[7]~5_combout ),
	.cout());
defparam \R_src2_lo[7]~5 .lut_mask = 16'hACFF;
defparam \R_src2_lo[7]~5 .sum_lutc_input = "datac";

dffeas \E_src2[7] (
	.clk(clk_clk),
	.d(\R_src2_lo[7]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[7]~q ),
	.prn(vcc));
defparam \E_src2[7] .is_wysiwyg = "true";
defparam \E_src2[7] .power_up = "low";

cycloneive_lcell_comb \Add1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[7]~q ),
	.cin(gnd),
	.combout(\Add1~5_combout ),
	.cout());
defparam \Add1~5 .lut_mask = 16'h0FF0;
defparam \Add1~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[7]~8 (
	.dataa(\D_iw[11]~q ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[7] ),
	.datac(gnd),
	.datad(\R_src1~36_combout ),
	.cin(gnd),
	.combout(\E_src1[7]~8_combout ),
	.cout());
defparam \E_src1[7]~8 .lut_mask = 16'hAACC;
defparam \E_src1[7]~8 .sum_lutc_input = "datac";

dffeas \E_src1[7] (
	.clk(clk_clk),
	.d(\E_src1[7]~8_combout ),
	.asdata(\F_pc_plus_one[5]~10_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~37_combout ),
	.ena(vcc),
	.q(\E_src1[7]~q ),
	.prn(vcc));
defparam \E_src1[7] .is_wysiwyg = "true";
defparam \E_src1[7] .power_up = "low";

cycloneive_lcell_comb \R_src2_lo[6]~6 (
	.dataa(\D_iw[12]~q ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[7]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[6]~6_combout ),
	.cout());
defparam \R_src2_lo[6]~6 .lut_mask = 16'hACFF;
defparam \R_src2_lo[6]~6 .sum_lutc_input = "datac";

dffeas \E_src2[6] (
	.clk(clk_clk),
	.d(\R_src2_lo[6]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[6]~q ),
	.prn(vcc));
defparam \E_src2[6] .is_wysiwyg = "true";
defparam \E_src2[6] .power_up = "low";

cycloneive_lcell_comb \Add1~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[6]~q ),
	.cin(gnd),
	.combout(\Add1~6_combout ),
	.cout());
defparam \Add1~6 .lut_mask = 16'h0FF0;
defparam \Add1~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[6]~9 (
	.dataa(\D_iw[10]~q ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[6] ),
	.datac(gnd),
	.datad(\R_src1~36_combout ),
	.cin(gnd),
	.combout(\E_src1[6]~9_combout ),
	.cout());
defparam \E_src1[6]~9 .lut_mask = 16'hAACC;
defparam \E_src1[6]~9 .sum_lutc_input = "datac";

dffeas \E_src1[6] (
	.clk(clk_clk),
	.d(\E_src1[6]~9_combout ),
	.asdata(\F_pc_plus_one[4]~8_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~37_combout ),
	.ena(vcc),
	.q(\E_src1[6]~q ),
	.prn(vcc));
defparam \E_src1[6] .is_wysiwyg = "true";
defparam \E_src1[6] .power_up = "low";

cycloneive_lcell_comb \R_src2_lo[5]~7 (
	.dataa(\D_iw[11]~q ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[7]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[5]~7_combout ),
	.cout());
defparam \R_src2_lo[5]~7 .lut_mask = 16'hACFF;
defparam \R_src2_lo[5]~7 .sum_lutc_input = "datac";

dffeas \E_src2[5] (
	.clk(clk_clk),
	.d(\R_src2_lo[5]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[5]~q ),
	.prn(vcc));
defparam \E_src2[5] .is_wysiwyg = "true";
defparam \E_src2[5] .power_up = "low";

cycloneive_lcell_comb \Add1~7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[5]~q ),
	.cin(gnd),
	.combout(\Add1~7_combout ),
	.cout());
defparam \Add1~7 .lut_mask = 16'h0FF0;
defparam \Add1~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[5]~10 (
	.dataa(\D_iw[9]~q ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[5] ),
	.datac(gnd),
	.datad(\R_src1~36_combout ),
	.cin(gnd),
	.combout(\E_src1[5]~10_combout ),
	.cout());
defparam \E_src1[5]~10 .lut_mask = 16'hAACC;
defparam \E_src1[5]~10 .sum_lutc_input = "datac";

dffeas \E_src1[5] (
	.clk(clk_clk),
	.d(\E_src1[5]~10_combout ),
	.asdata(\F_pc_plus_one[3]~6_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~37_combout ),
	.ena(vcc),
	.q(\E_src1[5]~q ),
	.prn(vcc));
defparam \E_src1[5] .is_wysiwyg = "true";
defparam \E_src1[5] .power_up = "low";

cycloneive_lcell_comb \Add1~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_src2[4]~q ),
	.datad(\E_alu_sub~q ),
	.cin(gnd),
	.combout(\Add1~8_combout ),
	.cout());
defparam \Add1~8 .lut_mask = 16'h0FF0;
defparam \Add1~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[4]~11 (
	.dataa(\D_iw[8]~q ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[4] ),
	.datac(gnd),
	.datad(\R_src1~36_combout ),
	.cin(gnd),
	.combout(\E_src1[4]~11_combout ),
	.cout());
defparam \E_src1[4]~11 .lut_mask = 16'hAACC;
defparam \E_src1[4]~11 .sum_lutc_input = "datac";

dffeas \E_src1[4] (
	.clk(clk_clk),
	.d(\E_src1[4]~11_combout ),
	.asdata(\F_pc_plus_one[2]~4_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~37_combout ),
	.ena(vcc),
	.q(\E_src1[4]~q ),
	.prn(vcc));
defparam \E_src1[4] .is_wysiwyg = "true";
defparam \E_src1[4] .power_up = "low";

cycloneive_lcell_comb \Add1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[3]~q ),
	.cin(gnd),
	.combout(\Add1~9_combout ),
	.cout());
defparam \Add1~9 .lut_mask = 16'h0FF0;
defparam \Add1~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[3]~12 (
	.dataa(\D_iw[7]~q ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[3] ),
	.datac(gnd),
	.datad(\R_src1~36_combout ),
	.cin(gnd),
	.combout(\E_src1[3]~12_combout ),
	.cout());
defparam \E_src1[3]~12 .lut_mask = 16'hAACC;
defparam \E_src1[3]~12 .sum_lutc_input = "datac";

dffeas \E_src1[3] (
	.clk(clk_clk),
	.d(\E_src1[3]~12_combout ),
	.asdata(\F_pc_plus_one[1]~2_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~37_combout ),
	.ena(vcc),
	.q(\E_src1[3]~q ),
	.prn(vcc));
defparam \E_src1[3] .is_wysiwyg = "true";
defparam \E_src1[3] .power_up = "low";

cycloneive_lcell_comb \Add1~10 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[2]~q ),
	.cin(gnd),
	.combout(\Add1~10_combout ),
	.cout());
defparam \Add1~10 .lut_mask = 16'h0FF0;
defparam \Add1~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[2]~13 (
	.dataa(\D_iw[6]~q ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[2] ),
	.datac(gnd),
	.datad(\R_src1~36_combout ),
	.cin(gnd),
	.combout(\E_src1[2]~13_combout ),
	.cout());
defparam \E_src1[2]~13 .lut_mask = 16'hAACC;
defparam \E_src1[2]~13 .sum_lutc_input = "datac";

dffeas \E_src1[2] (
	.clk(clk_clk),
	.d(\E_src1[2]~13_combout ),
	.asdata(\F_pc_plus_one[0]~0_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~37_combout ),
	.ena(vcc),
	.q(\E_src1[2]~q ),
	.prn(vcc));
defparam \E_src1[2] .is_wysiwyg = "true";
defparam \E_src1[2] .power_up = "low";

cycloneive_lcell_comb \Add1~11 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[1]~q ),
	.cin(gnd),
	.combout(\Add1~11_combout ),
	.cout());
defparam \Add1~11 .lut_mask = 16'h0FF0;
defparam \Add1~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src1[1]~38 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[1] ),
	.datad(\R_src1~37_combout ),
	.cin(gnd),
	.combout(\R_src1[1]~38_combout ),
	.cout());
defparam \R_src1[1]~38 .lut_mask = 16'hF7FF;
defparam \R_src1[1]~38 .sum_lutc_input = "datac";

dffeas \E_src1[1] (
	.clk(clk_clk),
	.d(\R_src1[1]~38_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[1]~q ),
	.prn(vcc));
defparam \E_src1[1] .is_wysiwyg = "true";
defparam \E_src1[1] .power_up = "low";

cycloneive_lcell_comb \Add1~12 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[0]~q ),
	.cin(gnd),
	.combout(\Add1~12_combout ),
	.cout());
defparam \Add1~12 .lut_mask = 16'h0FF0;
defparam \Add1~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~14 (
	.dataa(\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\Add1~14_cout ));
defparam \Add1~14 .lut_mask = 16'h00AA;
defparam \Add1~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~15 (
	.dataa(\Add1~12_combout ),
	.datab(\E_src1[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~14_cout ),
	.combout(\Add1~15_combout ),
	.cout(\Add1~16 ));
defparam \Add1~15 .lut_mask = 16'h967F;
defparam \Add1~15 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~17 (
	.dataa(\Add1~11_combout ),
	.datab(\E_src1[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~16 ),
	.combout(\Add1~17_combout ),
	.cout(\Add1~18 ));
defparam \Add1~17 .lut_mask = 16'h96EF;
defparam \Add1~17 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~19 (
	.dataa(\Add1~10_combout ),
	.datab(\E_src1[2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~18 ),
	.combout(\Add1~19_combout ),
	.cout(\Add1~20 ));
defparam \Add1~19 .lut_mask = 16'h967F;
defparam \Add1~19 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~21 (
	.dataa(\Add1~9_combout ),
	.datab(\E_src1[3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~20 ),
	.combout(\Add1~21_combout ),
	.cout(\Add1~22 ));
defparam \Add1~21 .lut_mask = 16'h96EF;
defparam \Add1~21 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~23 (
	.dataa(\Add1~8_combout ),
	.datab(\E_src1[4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~22 ),
	.combout(\Add1~23_combout ),
	.cout(\Add1~24 ));
defparam \Add1~23 .lut_mask = 16'h967F;
defparam \Add1~23 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~25 (
	.dataa(\Add1~7_combout ),
	.datab(\E_src1[5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~24 ),
	.combout(\Add1~25_combout ),
	.cout(\Add1~26 ));
defparam \Add1~25 .lut_mask = 16'h96EF;
defparam \Add1~25 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~27 (
	.dataa(\Add1~6_combout ),
	.datab(\E_src1[6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~26 ),
	.combout(\Add1~27_combout ),
	.cout(\Add1~28 ));
defparam \Add1~27 .lut_mask = 16'h967F;
defparam \Add1~27 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~29 (
	.dataa(\Add1~5_combout ),
	.datab(\E_src1[7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~28 ),
	.combout(\Add1~29_combout ),
	.cout(\Add1~30 ));
defparam \Add1~29 .lut_mask = 16'h96EF;
defparam \Add1~29 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~31 (
	.dataa(\Add1~4_combout ),
	.datab(\E_src1[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~30 ),
	.combout(\Add1~31_combout ),
	.cout(\Add1~32 ));
defparam \Add1~31 .lut_mask = 16'h967F;
defparam \Add1~31 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~33 (
	.dataa(\Add1~3_combout ),
	.datab(\E_src1[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~32 ),
	.combout(\Add1~33_combout ),
	.cout(\Add1~34 ));
defparam \Add1~33 .lut_mask = 16'h96EF;
defparam \Add1~33 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~35 (
	.dataa(\Add1~2_combout ),
	.datab(\E_src1[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~34 ),
	.combout(\Add1~35_combout ),
	.cout(\Add1~36 ));
defparam \Add1~35 .lut_mask = 16'h967F;
defparam \Add1~35 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~37 (
	.dataa(\Add1~1_combout ),
	.datab(\E_src1[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~36 ),
	.combout(\Add1~37_combout ),
	.cout(\Add1~38 ));
defparam \Add1~37 .lut_mask = 16'h96EF;
defparam \Add1~37 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~39 (
	.dataa(\Add1~0_combout ),
	.datab(\E_src1[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~38 ),
	.combout(\Add1~39_combout ),
	.cout(\Add1~40 ));
defparam \Add1~39 .lut_mask = 16'h967F;
defparam \Add1~39 .sum_lutc_input = "cin";

cycloneive_lcell_comb \D_logic_op_raw[1]~0 (
	.dataa(\D_iw[4]~q ),
	.datab(\D_iw[15]~q ),
	.datac(\Equal0~2_combout ),
	.datad(\D_iw[5]~q ),
	.cin(gnd),
	.combout(\D_logic_op_raw[1]~0_combout ),
	.cout());
defparam \D_logic_op_raw[1]~0 .lut_mask = 16'hEFFF;
defparam \D_logic_op_raw[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_alu_force_xor~10 (
	.dataa(\Equal62~0_combout ),
	.datab(\D_op_cmpge~0_combout ),
	.datac(\D_ctrl_alu_force_xor~14_combout ),
	.datad(\Equal0~3_combout ),
	.cin(gnd),
	.combout(\D_ctrl_alu_force_xor~10_combout ),
	.cout());
defparam \D_ctrl_alu_force_xor~10 .lut_mask = 16'hFEFF;
defparam \D_ctrl_alu_force_xor~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_alu_force_xor~11 (
	.dataa(\Equal0~5_combout ),
	.datab(\D_iw[5]~q ),
	.datac(\Equal0~4_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_alu_force_xor~11_combout ),
	.cout());
defparam \D_ctrl_alu_force_xor~11 .lut_mask = 16'hFEFF;
defparam \D_ctrl_alu_force_xor~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_alu_force_xor~13 (
	.dataa(\D_iw[15]~q ),
	.datab(\D_iw[14]~q ),
	.datac(\Equal62~0_combout ),
	.datad(\Equal62~1_combout ),
	.cin(gnd),
	.combout(\D_ctrl_alu_force_xor~13_combout ),
	.cout());
defparam \D_ctrl_alu_force_xor~13 .lut_mask = 16'hFFD8;
defparam \D_ctrl_alu_force_xor~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_alu_force_xor~12 (
	.dataa(\D_ctrl_alu_force_xor~10_combout ),
	.datab(\D_ctrl_alu_force_xor~11_combout ),
	.datac(\Equal0~7_combout ),
	.datad(\D_ctrl_alu_force_xor~13_combout ),
	.cin(gnd),
	.combout(\D_ctrl_alu_force_xor~12_combout ),
	.cout());
defparam \D_ctrl_alu_force_xor~12 .lut_mask = 16'hFFFE;
defparam \D_ctrl_alu_force_xor~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_logic_op[1]~0 (
	.dataa(\D_logic_op_raw[1]~0_combout ),
	.datab(\D_ctrl_alu_force_xor~12_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_logic_op[1]~0_combout ),
	.cout());
defparam \D_logic_op[1]~0 .lut_mask = 16'hEEEE;
defparam \D_logic_op[1]~0 .sum_lutc_input = "datac";

dffeas \R_logic_op[1] (
	.clk(clk_clk),
	.d(\D_logic_op[1]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_logic_op[1]~q ),
	.prn(vcc));
defparam \R_logic_op[1] .is_wysiwyg = "true";
defparam \R_logic_op[1] .power_up = "low";

cycloneive_lcell_comb \D_logic_op[0]~1 (
	.dataa(\D_ctrl_alu_force_xor~12_combout ),
	.datab(\D_iw[14]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\Equal0~7_combout ),
	.cin(gnd),
	.combout(\D_logic_op[0]~1_combout ),
	.cout());
defparam \D_logic_op[0]~1 .lut_mask = 16'hFAFC;
defparam \D_logic_op[0]~1 .sum_lutc_input = "datac";

dffeas \R_logic_op[0] (
	.clk(clk_clk),
	.d(\D_logic_op[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_logic_op[0]~q ),
	.prn(vcc));
defparam \R_logic_op[0] .is_wysiwyg = "true";
defparam \R_logic_op[0] .power_up = "low";

cycloneive_lcell_comb \E_logic_result[12]~0 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[12]~q ),
	.datac(\E_src1[12]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[12]~0_combout ),
	.cout());
defparam \E_logic_result[12]~0 .lut_mask = 16'h6996;
defparam \E_logic_result[12]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~8 (
	.dataa(\D_iw[13]~q ),
	.datab(gnd),
	.datac(\D_iw[11]~q ),
	.datad(\D_iw[16]~q ),
	.cin(gnd),
	.combout(\Equal0~8_combout ),
	.cout());
defparam \Equal0~8 .lut_mask = 16'hAFFF;
defparam \Equal0~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~10 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~10_combout ),
	.cout());
defparam \Equal0~10 .lut_mask = 16'hFFF7;
defparam \Equal0~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_logic~0 (
	.dataa(gnd),
	.datab(\D_iw[4]~q ),
	.datac(\Equal0~9_combout ),
	.datad(\Equal0~10_combout ),
	.cin(gnd),
	.combout(\D_ctrl_logic~0_combout ),
	.cout());
defparam \D_ctrl_logic~0 .lut_mask = 16'h3FFF;
defparam \D_ctrl_logic~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb D_ctrl_logic(
	.dataa(\Equal0~7_combout ),
	.datab(\D_iw[12]~q ),
	.datac(\Equal0~8_combout ),
	.datad(\D_ctrl_logic~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_logic~combout ),
	.cout());
defparam D_ctrl_logic.lut_mask = 16'hFEFF;
defparam D_ctrl_logic.sum_lutc_input = "datac";

dffeas R_ctrl_logic(
	.clk(clk_clk),
	.d(\D_ctrl_logic~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_logic~q ),
	.prn(vcc));
defparam R_ctrl_logic.is_wysiwyg = "true";
defparam R_ctrl_logic.power_up = "low";

cycloneive_lcell_comb \W_alu_result[12]~3 (
	.dataa(\Add1~39_combout ),
	.datab(\E_logic_result[12]~0_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[12]~3_combout ),
	.cout());
defparam \W_alu_result[12]~3 .lut_mask = 16'hAACC;
defparam \W_alu_result[12]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_shift_rot_right~0 (
	.dataa(\D_iw[11]~q ),
	.datab(\D_iw[12]~q ),
	.datac(\D_iw[15]~q ),
	.datad(\D_iw[16]~q ),
	.cin(gnd),
	.combout(\D_ctrl_shift_rot_right~0_combout ),
	.cout());
defparam \D_ctrl_shift_rot_right~0 .lut_mask = 16'hFEFF;
defparam \D_ctrl_shift_rot_right~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_shift_rot_right~1 (
	.dataa(\Equal0~7_combout ),
	.datab(\D_iw[14]~q ),
	.datac(\D_ctrl_shift_rot_right~0_combout ),
	.datad(\D_iw[13]~q ),
	.cin(gnd),
	.combout(\D_ctrl_shift_rot_right~1_combout ),
	.cout());
defparam \D_ctrl_shift_rot_right~1 .lut_mask = 16'hFEFF;
defparam \D_ctrl_shift_rot_right~1 .sum_lutc_input = "datac";

dffeas R_ctrl_shift_rot_right(
	.clk(clk_clk),
	.d(\D_ctrl_shift_rot_right~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_shift_rot_right~q ),
	.prn(vcc));
defparam R_ctrl_shift_rot_right.is_wysiwyg = "true";
defparam R_ctrl_shift_rot_right.power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[11]~4 (
	.dataa(\E_shift_rot_result[12]~q ),
	.datab(\E_shift_rot_result[10]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[11]~4_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[11]~4 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[11]~4 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[11] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[11]~4_combout ),
	.asdata(\E_src1[11]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[11]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[11] .is_wysiwyg = "true";
defparam \E_shift_rot_result[11] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[10]~5 (
	.dataa(\E_shift_rot_result[11]~q ),
	.datab(\E_shift_rot_result[9]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[10]~5_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[10]~5 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[10]~5 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[10] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[10]~5_combout ),
	.asdata(\E_src1[10]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[10]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[10] .is_wysiwyg = "true";
defparam \E_shift_rot_result[10] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[9]~6 (
	.dataa(\E_shift_rot_result[10]~q ),
	.datab(\E_shift_rot_result[8]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[9]~6_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[9]~6 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[9]~6 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[9] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[9]~6_combout ),
	.asdata(\E_src1[9]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[9]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[9] .is_wysiwyg = "true";
defparam \E_shift_rot_result[9] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[8]~7 (
	.dataa(\E_shift_rot_result[9]~q ),
	.datab(\E_shift_rot_result[7]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[8]~7_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[8]~7 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[8]~7 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[8] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[8]~7_combout ),
	.asdata(\E_src1[8]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[8]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[8] .is_wysiwyg = "true";
defparam \E_shift_rot_result[8] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[7]~8 (
	.dataa(\E_shift_rot_result[8]~q ),
	.datab(\E_shift_rot_result[6]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[7]~8_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[7]~8 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[7]~8 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[7] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[7]~8_combout ),
	.asdata(\E_src1[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[7]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[7] .is_wysiwyg = "true";
defparam \E_shift_rot_result[7] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[6]~9 (
	.dataa(\E_shift_rot_result[7]~q ),
	.datab(\E_shift_rot_result[5]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[6]~9_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[6]~9 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[6]~9 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[6] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[6]~9_combout ),
	.asdata(\E_src1[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[6]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[6] .is_wysiwyg = "true";
defparam \E_shift_rot_result[6] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[5]~10 (
	.dataa(\E_shift_rot_result[6]~q ),
	.datab(\E_shift_rot_result[4]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[5]~10_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[5]~10 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[5]~10 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[5] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[5]~10_combout ),
	.asdata(\E_src1[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[5]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[5] .is_wysiwyg = "true";
defparam \E_shift_rot_result[5] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[4]~11 (
	.dataa(\E_shift_rot_result[5]~q ),
	.datab(\E_shift_rot_result[3]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[4]~11_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[4]~11 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[4]~11 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[4] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[4]~11_combout ),
	.asdata(\E_src1[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[4]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[4] .is_wysiwyg = "true";
defparam \E_shift_rot_result[4] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[3]~12 (
	.dataa(\E_shift_rot_result[4]~q ),
	.datab(\E_shift_rot_result[2]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[3]~12_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[3]~12 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[3]~12 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[3] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[3]~12_combout ),
	.asdata(\E_src1[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[3]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[3] .is_wysiwyg = "true";
defparam \E_shift_rot_result[3] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[2]~13 (
	.dataa(\E_shift_rot_result[3]~q ),
	.datab(\E_shift_rot_result[1]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[2]~13_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[2]~13 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[2]~13 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[2] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[2]~13_combout ),
	.asdata(\E_src1[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[2]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[2] .is_wysiwyg = "true";
defparam \E_shift_rot_result[2] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[1]~15 (
	.dataa(\E_shift_rot_result[2]~q ),
	.datab(\E_shift_rot_result[0]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[1]~15_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[1]~15 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[1]~15 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[1] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[1]~15_combout ),
	.asdata(\E_src1[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[1]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[1] .is_wysiwyg = "true";
defparam \E_shift_rot_result[1] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[0]~16 (
	.dataa(\E_shift_rot_result[1]~q ),
	.datab(\E_shift_rot_fill_bit~0_combout ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[0]~16_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[0]~16 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[0]~16 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[0] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[0]~16_combout ),
	.asdata(\E_src1[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[0]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[0] .is_wysiwyg = "true";
defparam \E_shift_rot_result[0] .power_up = "low";

cycloneive_lcell_comb \R_ctrl_rot_right_nxt~0 (
	.dataa(\Equal0~7_combout ),
	.datab(\D_iw[14]~q ),
	.datac(\Equal62~7_combout ),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\R_ctrl_rot_right_nxt~0_combout ),
	.cout());
defparam \R_ctrl_rot_right_nxt~0 .lut_mask = 16'hFEFF;
defparam \R_ctrl_rot_right_nxt~0 .sum_lutc_input = "datac";

dffeas R_ctrl_rot_right(
	.clk(clk_clk),
	.d(\R_ctrl_rot_right_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_rot_right~q ),
	.prn(vcc));
defparam R_ctrl_rot_right.is_wysiwyg = "true";
defparam R_ctrl_rot_right.power_up = "low";

cycloneive_lcell_comb \D_ctrl_shift_logical~1 (
	.dataa(\D_ctrl_shift_logical~0_combout ),
	.datab(\D_iw[14]~q ),
	.datac(\Equal62~4_combout ),
	.datad(\Equal62~7_combout ),
	.cin(gnd),
	.combout(\D_ctrl_shift_logical~1_combout ),
	.cout());
defparam \D_ctrl_shift_logical~1 .lut_mask = 16'hFFB8;
defparam \D_ctrl_shift_logical~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_shift_logical~2 (
	.dataa(\Equal0~7_combout ),
	.datab(\D_iw[15]~q ),
	.datac(\D_ctrl_shift_logical~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_shift_logical~2_combout ),
	.cout());
defparam \D_ctrl_shift_logical~2 .lut_mask = 16'hFEFE;
defparam \D_ctrl_shift_logical~2 .sum_lutc_input = "datac";

dffeas R_ctrl_shift_logical(
	.clk(clk_clk),
	.d(\D_ctrl_shift_logical~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_shift_logical~q ),
	.prn(vcc));
defparam R_ctrl_shift_logical.is_wysiwyg = "true";
defparam R_ctrl_shift_logical.power_up = "low";

cycloneive_lcell_comb \E_shift_rot_fill_bit~0 (
	.dataa(\E_shift_rot_result[0]~q ),
	.datab(\E_shift_rot_result[31]~q ),
	.datac(\R_ctrl_rot_right~q ),
	.datad(\R_ctrl_shift_logical~q ),
	.cin(gnd),
	.combout(\E_shift_rot_fill_bit~0_combout ),
	.cout());
defparam \E_shift_rot_fill_bit~0 .lut_mask = 16'hACFF;
defparam \E_shift_rot_fill_bit~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_shift_rot_result_nxt[31]~18 (
	.dataa(\E_shift_rot_fill_bit~0_combout ),
	.datab(\E_shift_rot_result[30]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[31]~18_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[31]~18 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[31]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src1[31]~40 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[31] ),
	.datad(\R_src1~37_combout ),
	.cin(gnd),
	.combout(\R_src1[31]~40_combout ),
	.cout());
defparam \R_src1[31]~40 .lut_mask = 16'hF7FF;
defparam \R_src1[31]~40 .sum_lutc_input = "datac";

dffeas \E_src1[31] (
	.clk(clk_clk),
	.d(\R_src1[31]~40_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[31]~q ),
	.prn(vcc));
defparam \E_src1[31] .is_wysiwyg = "true";
defparam \E_src1[31] .power_up = "low";

dffeas \E_shift_rot_result[31] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[31]~18_combout ),
	.asdata(\E_src1[31]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[31]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[31] .is_wysiwyg = "true";
defparam \E_shift_rot_result[31] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[30]~20 (
	.dataa(\E_shift_rot_result[31]~q ),
	.datab(\E_shift_rot_result[29]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[30]~20_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[30]~20 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[30]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src1[30]~42 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[30] ),
	.datad(\R_src1~37_combout ),
	.cin(gnd),
	.combout(\R_src1[30]~42_combout ),
	.cout());
defparam \R_src1[30]~42 .lut_mask = 16'hF7FF;
defparam \R_src1[30]~42 .sum_lutc_input = "datac";

dffeas \E_src1[30] (
	.clk(clk_clk),
	.d(\R_src1[30]~42_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[30]~q ),
	.prn(vcc));
defparam \E_src1[30] .is_wysiwyg = "true";
defparam \E_src1[30] .power_up = "low";

dffeas \E_shift_rot_result[30] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[30]~20_combout ),
	.asdata(\E_src1[30]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[30]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[30] .is_wysiwyg = "true";
defparam \E_shift_rot_result[30] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[29]~22 (
	.dataa(\E_shift_rot_result[30]~q ),
	.datab(\E_shift_rot_result[28]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[29]~22_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[29]~22 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[29]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src1[29]~43 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[29] ),
	.datad(\R_src1~37_combout ),
	.cin(gnd),
	.combout(\R_src1[29]~43_combout ),
	.cout());
defparam \R_src1[29]~43 .lut_mask = 16'hF7FF;
defparam \R_src1[29]~43 .sum_lutc_input = "datac";

dffeas \E_src1[29] (
	.clk(clk_clk),
	.d(\R_src1[29]~43_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[29]~q ),
	.prn(vcc));
defparam \E_src1[29] .is_wysiwyg = "true";
defparam \E_src1[29] .power_up = "low";

dffeas \E_shift_rot_result[29] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[29]~22_combout ),
	.asdata(\E_src1[29]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[29]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[29] .is_wysiwyg = "true";
defparam \E_shift_rot_result[29] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[28]~23 (
	.dataa(\E_shift_rot_result[29]~q ),
	.datab(\E_shift_rot_result[27]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[28]~23_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[28]~23 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[28]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src1[28]~44 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[28] ),
	.datad(\R_src1~37_combout ),
	.cin(gnd),
	.combout(\R_src1[28]~44_combout ),
	.cout());
defparam \R_src1[28]~44 .lut_mask = 16'hF7FF;
defparam \R_src1[28]~44 .sum_lutc_input = "datac";

dffeas \E_src1[28] (
	.clk(clk_clk),
	.d(\R_src1[28]~44_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[28]~q ),
	.prn(vcc));
defparam \E_src1[28] .is_wysiwyg = "true";
defparam \E_src1[28] .power_up = "low";

dffeas \E_shift_rot_result[28] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[28]~23_combout ),
	.asdata(\E_src1[28]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[28]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[28] .is_wysiwyg = "true";
defparam \E_shift_rot_result[28] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[27]~24 (
	.dataa(\E_shift_rot_result[28]~q ),
	.datab(\E_shift_rot_result[26]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[27]~24_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[27]~24 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[27]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src1[27]~45 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[27] ),
	.datad(\R_src1~37_combout ),
	.cin(gnd),
	.combout(\R_src1[27]~45_combout ),
	.cout());
defparam \R_src1[27]~45 .lut_mask = 16'hF7FF;
defparam \R_src1[27]~45 .sum_lutc_input = "datac";

dffeas \E_src1[27] (
	.clk(clk_clk),
	.d(\R_src1[27]~45_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[27]~q ),
	.prn(vcc));
defparam \E_src1[27] .is_wysiwyg = "true";
defparam \E_src1[27] .power_up = "low";

dffeas \E_shift_rot_result[27] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[27]~24_combout ),
	.asdata(\E_src1[27]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[27]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[27] .is_wysiwyg = "true";
defparam \E_shift_rot_result[27] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[26]~25 (
	.dataa(\E_shift_rot_result[27]~q ),
	.datab(\E_shift_rot_result[25]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[26]~25_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[26]~25 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[26]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src1[26]~46 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[26] ),
	.datad(\R_src1~37_combout ),
	.cin(gnd),
	.combout(\R_src1[26]~46_combout ),
	.cout());
defparam \R_src1[26]~46 .lut_mask = 16'hF7FF;
defparam \R_src1[26]~46 .sum_lutc_input = "datac";

dffeas \E_src1[26] (
	.clk(clk_clk),
	.d(\R_src1[26]~46_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[26]~q ),
	.prn(vcc));
defparam \E_src1[26] .is_wysiwyg = "true";
defparam \E_src1[26] .power_up = "low";

dffeas \E_shift_rot_result[26] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[26]~25_combout ),
	.asdata(\E_src1[26]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[26]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[26] .is_wysiwyg = "true";
defparam \E_shift_rot_result[26] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[25]~26 (
	.dataa(\E_shift_rot_result[26]~q ),
	.datab(\E_shift_rot_result[24]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[25]~26_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[25]~26 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[25]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src1[25]~47 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[25] ),
	.datad(\R_src1~37_combout ),
	.cin(gnd),
	.combout(\R_src1[25]~47_combout ),
	.cout());
defparam \R_src1[25]~47 .lut_mask = 16'hF7FF;
defparam \R_src1[25]~47 .sum_lutc_input = "datac";

dffeas \E_src1[25] (
	.clk(clk_clk),
	.d(\R_src1[25]~47_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[25]~q ),
	.prn(vcc));
defparam \E_src1[25] .is_wysiwyg = "true";
defparam \E_src1[25] .power_up = "low";

dffeas \E_shift_rot_result[25] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[25]~26_combout ),
	.asdata(\E_src1[25]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[25]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[25] .is_wysiwyg = "true";
defparam \E_shift_rot_result[25] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[24]~27 (
	.dataa(\E_shift_rot_result[25]~q ),
	.datab(\E_shift_rot_result[23]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[24]~27_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[24]~27 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[24]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src1[24]~48 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[24] ),
	.datad(\R_src1~37_combout ),
	.cin(gnd),
	.combout(\R_src1[24]~48_combout ),
	.cout());
defparam \R_src1[24]~48 .lut_mask = 16'hF7FF;
defparam \R_src1[24]~48 .sum_lutc_input = "datac";

dffeas \E_src1[24] (
	.clk(clk_clk),
	.d(\R_src1[24]~48_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[24]~q ),
	.prn(vcc));
defparam \E_src1[24] .is_wysiwyg = "true";
defparam \E_src1[24] .power_up = "low";

dffeas \E_shift_rot_result[24] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[24]~27_combout ),
	.asdata(\E_src1[24]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[24]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[24] .is_wysiwyg = "true";
defparam \E_shift_rot_result[24] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[23]~28 (
	.dataa(\E_shift_rot_result[24]~q ),
	.datab(\E_shift_rot_result[22]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[23]~28_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[23]~28 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[23]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src1[23]~49 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[23] ),
	.datad(\R_src1~37_combout ),
	.cin(gnd),
	.combout(\R_src1[23]~49_combout ),
	.cout());
defparam \R_src1[23]~49 .lut_mask = 16'hF7FF;
defparam \R_src1[23]~49 .sum_lutc_input = "datac";

dffeas \E_src1[23] (
	.clk(clk_clk),
	.d(\R_src1[23]~49_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[23]~q ),
	.prn(vcc));
defparam \E_src1[23] .is_wysiwyg = "true";
defparam \E_src1[23] .power_up = "low";

dffeas \E_shift_rot_result[23] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[23]~28_combout ),
	.asdata(\E_src1[23]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[23]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[23] .is_wysiwyg = "true";
defparam \E_shift_rot_result[23] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[22]~29 (
	.dataa(\E_shift_rot_result[23]~q ),
	.datab(\E_shift_rot_result[21]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[22]~29_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[22]~29 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[22]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src1[22]~50 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[22] ),
	.datad(\R_src1~37_combout ),
	.cin(gnd),
	.combout(\R_src1[22]~50_combout ),
	.cout());
defparam \R_src1[22]~50 .lut_mask = 16'hF7FF;
defparam \R_src1[22]~50 .sum_lutc_input = "datac";

dffeas \E_src1[22] (
	.clk(clk_clk),
	.d(\R_src1[22]~50_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[22]~q ),
	.prn(vcc));
defparam \E_src1[22] .is_wysiwyg = "true";
defparam \E_src1[22] .power_up = "low";

dffeas \E_shift_rot_result[22] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[22]~29_combout ),
	.asdata(\E_src1[22]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[22]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[22] .is_wysiwyg = "true";
defparam \E_shift_rot_result[22] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[21]~30 (
	.dataa(\E_shift_rot_result[22]~q ),
	.datab(\E_shift_rot_result[20]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[21]~30_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[21]~30 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[21]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src1[21]~51 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[21] ),
	.datad(\R_src1~37_combout ),
	.cin(gnd),
	.combout(\R_src1[21]~51_combout ),
	.cout());
defparam \R_src1[21]~51 .lut_mask = 16'hF7FF;
defparam \R_src1[21]~51 .sum_lutc_input = "datac";

dffeas \E_src1[21] (
	.clk(clk_clk),
	.d(\R_src1[21]~51_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[21]~q ),
	.prn(vcc));
defparam \E_src1[21] .is_wysiwyg = "true";
defparam \E_src1[21] .power_up = "low";

dffeas \E_shift_rot_result[21] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[21]~30_combout ),
	.asdata(\E_src1[21]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[21]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[21] .is_wysiwyg = "true";
defparam \E_shift_rot_result[21] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[20]~31 (
	.dataa(\E_shift_rot_result[21]~q ),
	.datab(\E_shift_rot_result[19]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[20]~31_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[20]~31 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[20]~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src1[20]~52 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[20] ),
	.datad(\R_src1~37_combout ),
	.cin(gnd),
	.combout(\R_src1[20]~52_combout ),
	.cout());
defparam \R_src1[20]~52 .lut_mask = 16'hF7FF;
defparam \R_src1[20]~52 .sum_lutc_input = "datac";

dffeas \E_src1[20] (
	.clk(clk_clk),
	.d(\R_src1[20]~52_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[20]~q ),
	.prn(vcc));
defparam \E_src1[20] .is_wysiwyg = "true";
defparam \E_src1[20] .power_up = "low";

dffeas \E_shift_rot_result[20] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[20]~31_combout ),
	.asdata(\E_src1[20]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[20]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[20] .is_wysiwyg = "true";
defparam \E_shift_rot_result[20] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[19]~21 (
	.dataa(\E_shift_rot_result[20]~q ),
	.datab(\E_shift_rot_result[18]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[19]~21_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[19]~21 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[19]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src1[19]~53 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[19] ),
	.datad(\R_src1~37_combout ),
	.cin(gnd),
	.combout(\R_src1[19]~53_combout ),
	.cout());
defparam \R_src1[19]~53 .lut_mask = 16'hF7FF;
defparam \R_src1[19]~53 .sum_lutc_input = "datac";

dffeas \E_src1[19] (
	.clk(clk_clk),
	.d(\R_src1[19]~53_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[19]~q ),
	.prn(vcc));
defparam \E_src1[19] .is_wysiwyg = "true";
defparam \E_src1[19] .power_up = "low";

dffeas \E_shift_rot_result[19] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[19]~21_combout ),
	.asdata(\E_src1[19]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[19]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[19] .is_wysiwyg = "true";
defparam \E_shift_rot_result[19] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[18]~19 (
	.dataa(\E_shift_rot_result[19]~q ),
	.datab(\E_shift_rot_result[17]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[18]~19_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[18]~19 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[18]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src1[18]~54 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[18] ),
	.datad(\R_src1~37_combout ),
	.cin(gnd),
	.combout(\R_src1[18]~54_combout ),
	.cout());
defparam \R_src1[18]~54 .lut_mask = 16'hF7FF;
defparam \R_src1[18]~54 .sum_lutc_input = "datac";

dffeas \E_src1[18] (
	.clk(clk_clk),
	.d(\R_src1[18]~54_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[18]~q ),
	.prn(vcc));
defparam \E_src1[18] .is_wysiwyg = "true";
defparam \E_src1[18] .power_up = "low";

dffeas \E_shift_rot_result[18] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[18]~19_combout ),
	.asdata(\E_src1[18]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[18]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[18] .is_wysiwyg = "true";
defparam \E_shift_rot_result[18] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[17]~17 (
	.dataa(\E_shift_rot_result[18]~q ),
	.datab(\E_shift_rot_result[16]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[17]~17_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[17]~17 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[17]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src1[17]~55 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[17] ),
	.datad(\R_src1~37_combout ),
	.cin(gnd),
	.combout(\R_src1[17]~55_combout ),
	.cout());
defparam \R_src1[17]~55 .lut_mask = 16'hF7FF;
defparam \R_src1[17]~55 .sum_lutc_input = "datac";

dffeas \E_src1[17] (
	.clk(clk_clk),
	.d(\R_src1[17]~55_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[17]~q ),
	.prn(vcc));
defparam \E_src1[17] .is_wysiwyg = "true";
defparam \E_src1[17] .power_up = "low";

dffeas \E_shift_rot_result[17] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[17]~17_combout ),
	.asdata(\E_src1[17]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[17]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[17] .is_wysiwyg = "true";
defparam \E_shift_rot_result[17] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[16]~14 (
	.dataa(\E_shift_rot_result[17]~q ),
	.datab(\E_shift_rot_result[15]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[16]~14_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[16]~14 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[16]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src1[16]~41 (
	.dataa(\E_valid_from_R~q ),
	.datab(\R_ctrl_jmp_direct~q ),
	.datac(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[16] ),
	.datad(\R_src1~37_combout ),
	.cin(gnd),
	.combout(\R_src1[16]~41_combout ),
	.cout());
defparam \R_src1[16]~41 .lut_mask = 16'hF7FF;
defparam \R_src1[16]~41 .sum_lutc_input = "datac";

dffeas \E_src1[16] (
	.clk(clk_clk),
	.d(\R_src1[16]~41_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src1[16]~q ),
	.prn(vcc));
defparam \E_src1[16] .is_wysiwyg = "true";
defparam \E_src1[16] .power_up = "low";

dffeas \E_shift_rot_result[16] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[16]~14_combout ),
	.asdata(\E_src1[16]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[16]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[16] .is_wysiwyg = "true";
defparam \E_shift_rot_result[16] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[15]~1 (
	.dataa(\E_shift_rot_result[16]~q ),
	.datab(\E_shift_rot_result[14]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[15]~1_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[15]~1 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[15]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[19]~41 (
	.dataa(src_payload9),
	.datab(src1_valid),
	.datac(av_readdata_pre_19),
	.datad(\D_iw[27]~0_combout ),
	.cin(gnd),
	.combout(\F_iw[19]~41_combout ),
	.cout());
defparam \F_iw[19]~41 .lut_mask = 16'hFEFF;
defparam \F_iw[19]~41 .sum_lutc_input = "datac";

dffeas \D_iw[19] (
	.clk(clk_clk),
	.d(\F_iw[19]~41_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[19]~q ),
	.prn(vcc));
defparam \D_iw[19] .is_wysiwyg = "true";
defparam \D_iw[19] .power_up = "low";

cycloneive_lcell_comb \E_src1[15]~0 (
	.dataa(\D_iw[19]~q ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[15] ),
	.datac(gnd),
	.datad(\R_src1~36_combout ),
	.cin(gnd),
	.combout(\E_src1[15]~0_combout ),
	.cout());
defparam \E_src1[15]~0 .lut_mask = 16'hAACC;
defparam \E_src1[15]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_plus_one[11]~22 (
	.dataa(F_pc_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[10]~21 ),
	.combout(\F_pc_plus_one[11]~22_combout ),
	.cout(\F_pc_plus_one[11]~23 ));
defparam \F_pc_plus_one[11]~22 .lut_mask = 16'h5A5F;
defparam \F_pc_plus_one[11]~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[12]~24 (
	.dataa(F_pc_12),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\F_pc_plus_one[11]~23 ),
	.combout(\F_pc_plus_one[12]~24_combout ),
	.cout(\F_pc_plus_one[12]~25 ));
defparam \F_pc_plus_one[12]~24 .lut_mask = 16'h5AAF;
defparam \F_pc_plus_one[12]~24 .sum_lutc_input = "cin";

cycloneive_lcell_comb \F_pc_plus_one[13]~26 (
	.dataa(F_pc_13),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\F_pc_plus_one[12]~25 ),
	.combout(\F_pc_plus_one[13]~26_combout ),
	.cout());
defparam \F_pc_plus_one[13]~26 .lut_mask = 16'h5A5A;
defparam \F_pc_plus_one[13]~26 .sum_lutc_input = "cin";

dffeas \E_src1[15] (
	.clk(clk_clk),
	.d(\E_src1[15]~0_combout ),
	.asdata(\F_pc_plus_one[13]~26_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~37_combout ),
	.ena(vcc),
	.q(\E_src1[15]~q ),
	.prn(vcc));
defparam \E_src1[15] .is_wysiwyg = "true";
defparam \E_src1[15] .power_up = "low";

dffeas \E_shift_rot_result[15] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[15]~1_combout ),
	.asdata(\E_src1[15]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[15]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[15] .is_wysiwyg = "true";
defparam \E_shift_rot_result[15] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[14]~2 (
	.dataa(\E_shift_rot_result[15]~q ),
	.datab(\E_shift_rot_result[13]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[14]~2_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[14]~2 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[14]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[14]~1 (
	.dataa(\D_iw[18]~q ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[14] ),
	.datac(gnd),
	.datad(\R_src1~36_combout ),
	.cin(gnd),
	.combout(\E_src1[14]~1_combout ),
	.cout());
defparam \E_src1[14]~1 .lut_mask = 16'hAACC;
defparam \E_src1[14]~1 .sum_lutc_input = "datac";

dffeas \E_src1[14] (
	.clk(clk_clk),
	.d(\E_src1[14]~1_combout ),
	.asdata(\F_pc_plus_one[12]~24_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~37_combout ),
	.ena(vcc),
	.q(\E_src1[14]~q ),
	.prn(vcc));
defparam \E_src1[14] .is_wysiwyg = "true";
defparam \E_src1[14] .power_up = "low";

dffeas \E_shift_rot_result[14] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[14]~2_combout ),
	.asdata(\E_src1[14]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[14]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[14] .is_wysiwyg = "true";
defparam \E_shift_rot_result[14] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[13]~3 (
	.dataa(\E_shift_rot_result[14]~q ),
	.datab(\E_shift_rot_result[12]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[13]~3_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[13]~3 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[13]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src1[13]~2 (
	.dataa(\D_iw[17]~q ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[13] ),
	.datac(gnd),
	.datad(\R_src1~36_combout ),
	.cin(gnd),
	.combout(\E_src1[13]~2_combout ),
	.cout());
defparam \E_src1[13]~2 .lut_mask = 16'hAACC;
defparam \E_src1[13]~2 .sum_lutc_input = "datac";

dffeas \E_src1[13] (
	.clk(clk_clk),
	.d(\E_src1[13]~2_combout ),
	.asdata(\F_pc_plus_one[11]~22_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\R_src1~37_combout ),
	.ena(vcc),
	.q(\E_src1[13]~q ),
	.prn(vcc));
defparam \E_src1[13] .is_wysiwyg = "true";
defparam \E_src1[13] .power_up = "low";

dffeas \E_shift_rot_result[13] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[13]~3_combout ),
	.asdata(\E_src1[13]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[13]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[13] .is_wysiwyg = "true";
defparam \E_shift_rot_result[13] .power_up = "low";

cycloneive_lcell_comb \E_shift_rot_result_nxt[12]~0 (
	.dataa(\E_shift_rot_result[13]~q ),
	.datab(\E_shift_rot_result[11]~q ),
	.datac(gnd),
	.datad(\R_ctrl_shift_rot_right~q ),
	.cin(gnd),
	.combout(\E_shift_rot_result_nxt[12]~0_combout ),
	.cout());
defparam \E_shift_rot_result_nxt[12]~0 .lut_mask = 16'hAACC;
defparam \E_shift_rot_result_nxt[12]~0 .sum_lutc_input = "datac";

dffeas \E_shift_rot_result[12] (
	.clk(clk_clk),
	.d(\E_shift_rot_result_nxt[12]~0_combout ),
	.asdata(\E_src1[12]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_new_inst~q ),
	.ena(vcc),
	.q(\E_shift_rot_result[12]~q ),
	.prn(vcc));
defparam \E_shift_rot_result[12] .is_wysiwyg = "true";
defparam \E_shift_rot_result[12] .power_up = "low";

cycloneive_lcell_comb D_op_rdctl(
	.dataa(\Equal0~7_combout ),
	.datab(\Equal62~3_combout ),
	.datac(\D_iw[15]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\D_op_rdctl~combout ),
	.cout());
defparam D_op_rdctl.lut_mask = 16'hEFFF;
defparam D_op_rdctl.sum_lutc_input = "datac";

dffeas R_ctrl_rd_ctl_reg(
	.clk(clk_clk),
	.d(\D_op_rdctl~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_rd_ctl_reg~q ),
	.prn(vcc));
defparam R_ctrl_rd_ctl_reg.is_wysiwyg = "true";
defparam R_ctrl_rd_ctl_reg.power_up = "low";

cycloneive_lcell_comb \Equal0~6 (
	.dataa(\D_iw[1]~q ),
	.datab(\D_iw[0]~q ),
	.datac(\D_iw[3]~q ),
	.datad(\D_iw[2]~q ),
	.cin(gnd),
	.combout(\Equal0~6_combout ),
	.cout());
defparam \Equal0~6 .lut_mask = 16'hF7FF;
defparam \Equal0~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_br_cmp~2 (
	.dataa(\Equal0~6_combout ),
	.datab(\Equal0~4_combout ),
	.datac(\Equal0~3_combout ),
	.datad(\D_ctrl_jmp_direct~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_br_cmp~2_combout ),
	.cout());
defparam \D_ctrl_br_cmp~2 .lut_mask = 16'hEFFF;
defparam \D_ctrl_br_cmp~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_br_cmp~5 (
	.dataa(\D_iw[15]~q ),
	.datab(\D_iw[14]~q ),
	.datac(\Equal62~0_combout ),
	.datad(\Equal62~1_combout ),
	.cin(gnd),
	.combout(\D_ctrl_br_cmp~5_combout ),
	.cout());
defparam \D_ctrl_br_cmp~5 .lut_mask = 16'hF7B3;
defparam \D_ctrl_br_cmp~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_br_cmp~3 (
	.dataa(\R_ctrl_br_nxt~1_combout ),
	.datab(\Equal0~7_combout ),
	.datac(\D_ctrl_br_cmp~5_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\D_ctrl_br_cmp~3_combout ),
	.cout());
defparam \D_ctrl_br_cmp~3 .lut_mask = 16'hFEFE;
defparam \D_ctrl_br_cmp~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_br_cmp~4 (
	.dataa(\D_ctrl_br_cmp~2_combout ),
	.datab(\D_ctrl_br_cmp~3_combout ),
	.datac(\Equal62~0_combout ),
	.datad(\D_op_cmpge~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_br_cmp~4_combout ),
	.cout());
defparam \D_ctrl_br_cmp~4 .lut_mask = 16'hFFFE;
defparam \D_ctrl_br_cmp~4 .sum_lutc_input = "datac";

dffeas R_ctrl_br_cmp(
	.clk(clk_clk),
	.d(\D_ctrl_br_cmp~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_br_cmp~q ),
	.prn(vcc));
defparam R_ctrl_br_cmp.is_wysiwyg = "true";
defparam R_ctrl_br_cmp.power_up = "low";

cycloneive_lcell_comb \E_alu_result~0 (
	.dataa(\R_ctrl_rd_ctl_reg~q ),
	.datab(\R_ctrl_br_cmp~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\E_alu_result~0_combout ),
	.cout());
defparam \E_alu_result~0 .lut_mask = 16'hEEEE;
defparam \E_alu_result~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[21]~40 (
	.dataa(src_payload8),
	.datab(src1_valid),
	.datac(av_readdata_pre_21),
	.datad(\D_iw[27]~0_combout ),
	.cin(gnd),
	.combout(\F_iw[21]~40_combout ),
	.cout());
defparam \F_iw[21]~40 .lut_mask = 16'hFEFF;
defparam \F_iw[21]~40 .sum_lutc_input = "datac";

dffeas \D_iw[21] (
	.clk(clk_clk),
	.d(\F_iw[21]~40_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[21]~q ),
	.prn(vcc));
defparam \D_iw[21] .is_wysiwyg = "true";
defparam \D_iw[21] .power_up = "low";

cycloneive_lcell_comb \R_src2_lo[15]~15 (
	.dataa(\D_iw[21]~q ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[7]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[15]~15_combout ),
	.cout());
defparam \R_src2_lo[15]~15 .lut_mask = 16'hACFF;
defparam \R_src2_lo[15]~15 .sum_lutc_input = "datac";

dffeas \E_src2[15] (
	.clk(clk_clk),
	.d(\R_src2_lo[15]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[15]~q ),
	.prn(vcc));
defparam \E_src2[15] .is_wysiwyg = "true";
defparam \E_src2[15] .power_up = "low";

cycloneive_lcell_comb \Add1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[15]~q ),
	.cin(gnd),
	.combout(\Add1~41_combout ),
	.cout());
defparam \Add1~41 .lut_mask = 16'h0FF0;
defparam \Add1~41 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_iw[20]~42 (
	.dataa(src_payload10),
	.datab(src1_valid),
	.datac(av_readdata_pre_20),
	.datad(\D_iw[27]~0_combout ),
	.cin(gnd),
	.combout(\F_iw[20]~42_combout ),
	.cout());
defparam \F_iw[20]~42 .lut_mask = 16'hFEFF;
defparam \F_iw[20]~42 .sum_lutc_input = "datac";

dffeas \D_iw[20] (
	.clk(clk_clk),
	.d(\F_iw[20]~42_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\F_valid~0_combout ),
	.q(\D_iw[20]~q ),
	.prn(vcc));
defparam \D_iw[20] .is_wysiwyg = "true";
defparam \D_iw[20] .power_up = "low";

cycloneive_lcell_comb \R_src2_lo[14]~16 (
	.dataa(\D_iw[20]~q ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[7]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[14]~16_combout ),
	.cout());
defparam \R_src2_lo[14]~16 .lut_mask = 16'hACFF;
defparam \R_src2_lo[14]~16 .sum_lutc_input = "datac";

dffeas \E_src2[14] (
	.clk(clk_clk),
	.d(\R_src2_lo[14]~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[14]~q ),
	.prn(vcc));
defparam \E_src2[14] .is_wysiwyg = "true";
defparam \E_src2[14] .power_up = "low";

cycloneive_lcell_comb \Add1~42 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[14]~q ),
	.cin(gnd),
	.combout(\Add1~42_combout ),
	.cout());
defparam \Add1~42 .lut_mask = 16'h0FF0;
defparam \Add1~42 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_lo[13]~17 (
	.dataa(\D_iw[19]~q ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\E_src2[7]~15_combout ),
	.cin(gnd),
	.combout(\R_src2_lo[13]~17_combout ),
	.cout());
defparam \R_src2_lo[13]~17 .lut_mask = 16'hACFF;
defparam \R_src2_lo[13]~17 .sum_lutc_input = "datac";

dffeas \E_src2[13] (
	.clk(clk_clk),
	.d(\R_src2_lo[13]~17_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[13]~q ),
	.prn(vcc));
defparam \E_src2[13] .is_wysiwyg = "true";
defparam \E_src2[13] .power_up = "low";

cycloneive_lcell_comb \Add1~43 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[13]~q ),
	.cin(gnd),
	.combout(\Add1~43_combout ),
	.cout());
defparam \Add1~43 .lut_mask = 16'h0FF0;
defparam \Add1~43 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~44 (
	.dataa(\Add1~43_combout ),
	.datab(\E_src1[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~40 ),
	.combout(\Add1~44_combout ),
	.cout(\Add1~45 ));
defparam \Add1~44 .lut_mask = 16'h96EF;
defparam \Add1~44 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~46 (
	.dataa(\Add1~42_combout ),
	.datab(\E_src1[14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~45 ),
	.combout(\Add1~46_combout ),
	.cout(\Add1~47 ));
defparam \Add1~46 .lut_mask = 16'h967F;
defparam \Add1~46 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add1~48 (
	.dataa(\Add1~41_combout ),
	.datab(\E_src1[15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~47 ),
	.combout(\Add1~48_combout ),
	.cout(\Add1~49 ));
defparam \Add1~48 .lut_mask = 16'h96EF;
defparam \Add1~48 .sum_lutc_input = "cin";

cycloneive_lcell_comb \E_logic_result[15]~1 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[15]~q ),
	.datac(\E_src1[15]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[15]~1_combout ),
	.cout());
defparam \E_logic_result[15]~1 .lut_mask = 16'h6996;
defparam \E_logic_result[15]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[15]~0 (
	.dataa(\Add1~48_combout ),
	.datab(\E_logic_result[15]~1_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[15]~0_combout ),
	.cout());
defparam \W_alu_result[15]~0 .lut_mask = 16'hAACC;
defparam \W_alu_result[15]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[14]~2 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[14]~q ),
	.datac(\E_src1[14]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[14]~2_combout ),
	.cout());
defparam \E_logic_result[14]~2 .lut_mask = 16'h6996;
defparam \E_logic_result[14]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[14]~1 (
	.dataa(\Add1~46_combout ),
	.datab(\E_logic_result[14]~2_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[14]~1_combout ),
	.cout());
defparam \W_alu_result[14]~1 .lut_mask = 16'hAACC;
defparam \W_alu_result[14]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[13]~3 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[13]~q ),
	.datac(\E_src1[13]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[13]~3_combout ),
	.cout());
defparam \E_logic_result[13]~3 .lut_mask = 16'h6996;
defparam \E_logic_result[13]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[13]~2 (
	.dataa(\Add1~44_combout ),
	.datab(\E_logic_result[13]~3_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[13]~2_combout ),
	.cout());
defparam \W_alu_result[13]~2 .lut_mask = 16'hAACC;
defparam \W_alu_result[13]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[11]~4 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[11]~q ),
	.datac(\E_src1[11]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[11]~4_combout ),
	.cout());
defparam \E_logic_result[11]~4 .lut_mask = 16'h6996;
defparam \E_logic_result[11]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[11]~4 (
	.dataa(\Add1~37_combout ),
	.datab(\E_logic_result[11]~4_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[11]~4_combout ),
	.cout());
defparam \W_alu_result[11]~4 .lut_mask = 16'hAACC;
defparam \W_alu_result[11]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[10]~5 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[10]~q ),
	.datac(\E_src1[10]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[10]~5_combout ),
	.cout());
defparam \E_logic_result[10]~5 .lut_mask = 16'h6996;
defparam \E_logic_result[10]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[10]~5 (
	.dataa(\Add1~35_combout ),
	.datab(\E_logic_result[10]~5_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[10]~5_combout ),
	.cout());
defparam \W_alu_result[10]~5 .lut_mask = 16'hAACC;
defparam \W_alu_result[10]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[9]~6 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[9]~q ),
	.datac(\E_src1[9]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[9]~6_combout ),
	.cout());
defparam \E_logic_result[9]~6 .lut_mask = 16'h6996;
defparam \E_logic_result[9]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[9]~6 (
	.dataa(\Add1~33_combout ),
	.datab(\E_logic_result[9]~6_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[9]~6_combout ),
	.cout());
defparam \W_alu_result[9]~6 .lut_mask = 16'hAACC;
defparam \W_alu_result[9]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[8]~7 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[8]~q ),
	.datac(\E_src1[8]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[8]~7_combout ),
	.cout());
defparam \E_logic_result[8]~7 .lut_mask = 16'h6996;
defparam \E_logic_result[8]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[8]~7 (
	.dataa(\Add1~31_combout ),
	.datab(\E_logic_result[8]~7_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[8]~7_combout ),
	.cout());
defparam \W_alu_result[8]~7 .lut_mask = 16'hAACC;
defparam \W_alu_result[8]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[7]~8 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[7]~q ),
	.datac(\E_src1[7]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[7]~8_combout ),
	.cout());
defparam \E_logic_result[7]~8 .lut_mask = 16'h6996;
defparam \E_logic_result[7]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[7]~8 (
	.dataa(\Add1~29_combout ),
	.datab(\E_logic_result[7]~8_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[7]~8_combout ),
	.cout());
defparam \W_alu_result[7]~8 .lut_mask = 16'hAACC;
defparam \W_alu_result[7]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[6]~9 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[6]~q ),
	.datac(\E_src1[6]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[6]~9_combout ),
	.cout());
defparam \E_logic_result[6]~9 .lut_mask = 16'h6996;
defparam \E_logic_result[6]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[6]~9 (
	.dataa(\Add1~27_combout ),
	.datab(\E_logic_result[6]~9_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[6]~9_combout ),
	.cout());
defparam \W_alu_result[6]~9 .lut_mask = 16'hAACC;
defparam \W_alu_result[6]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[5]~10 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[5]~q ),
	.datac(\E_src1[5]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[5]~10_combout ),
	.cout());
defparam \E_logic_result[5]~10 .lut_mask = 16'h6996;
defparam \E_logic_result[5]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[5]~10 (
	.dataa(\Add1~25_combout ),
	.datab(\E_logic_result[5]~10_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[5]~10_combout ),
	.cout());
defparam \W_alu_result[5]~10 .lut_mask = 16'hAACC;
defparam \W_alu_result[5]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[4]~11 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[4]~q ),
	.datac(\E_src1[4]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[4]~11_combout ),
	.cout());
defparam \E_logic_result[4]~11 .lut_mask = 16'h6996;
defparam \E_logic_result[4]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[4]~11 (
	.dataa(\Add1~23_combout ),
	.datab(\E_logic_result[4]~11_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[4]~11_combout ),
	.cout());
defparam \W_alu_result[4]~11 .lut_mask = 16'hAACC;
defparam \W_alu_result[4]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[3]~12 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[3]~q ),
	.datac(\E_src1[3]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[3]~12_combout ),
	.cout());
defparam \E_logic_result[3]~12 .lut_mask = 16'h6996;
defparam \E_logic_result[3]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[3]~12 (
	.dataa(\Add1~21_combout ),
	.datab(\E_logic_result[3]~12_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[3]~12_combout ),
	.cout());
defparam \W_alu_result[3]~12 .lut_mask = 16'hAACC;
defparam \W_alu_result[3]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[2]~13 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[2]~q ),
	.datac(\E_src1[2]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[2]~13_combout ),
	.cout());
defparam \E_logic_result[2]~13 .lut_mask = 16'h6996;
defparam \E_logic_result[2]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \W_alu_result[2]~13 (
	.dataa(\Add1~19_combout ),
	.datab(\E_logic_result[2]~13_combout ),
	.datac(gnd),
	.datad(\R_ctrl_logic~q ),
	.cin(gnd),
	.combout(\W_alu_result[2]~13_combout ),
	.cout());
defparam \W_alu_result[2]~13 .lut_mask = 16'hAACC;
defparam \W_alu_result[2]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \d_writedata[24]~0 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[24] ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[24]~0_combout ),
	.cout());
defparam \d_writedata[24]~0 .lut_mask = 16'hAACC;
defparam \d_writedata[24]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_mem8~0 (
	.dataa(\D_iw[0]~q ),
	.datab(\D_iw[1]~q ),
	.datac(\D_iw[2]~q ),
	.datad(\D_iw[3]~q ),
	.cin(gnd),
	.combout(\D_ctrl_mem8~0_combout ),
	.cout());
defparam \D_ctrl_mem8~0 .lut_mask = 16'hFEFF;
defparam \D_ctrl_mem8~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_mem8~1 (
	.dataa(\D_ctrl_mem8~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_mem8~1_combout ),
	.cout());
defparam \D_ctrl_mem8~1 .lut_mask = 16'hAAFF;
defparam \D_ctrl_mem8~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \d_writedata[25]~1 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[25] ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[25]~1_combout ),
	.cout());
defparam \d_writedata[25]~1 .lut_mask = 16'hAACC;
defparam \d_writedata[25]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \d_writedata[26]~2 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[26] ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[26]~2_combout ),
	.cout());
defparam \d_writedata[26]~2 .lut_mask = 16'hAACC;
defparam \d_writedata[26]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \d_writedata[27]~3 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[27] ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[27]~3_combout ),
	.cout());
defparam \d_writedata[27]~3 .lut_mask = 16'hAACC;
defparam \d_writedata[27]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \d_writedata[28]~4 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[28] ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[28]~4_combout ),
	.cout());
defparam \d_writedata[28]~4 .lut_mask = 16'hAACC;
defparam \d_writedata[28]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \d_writedata[29]~5 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[29] ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[29]~5_combout ),
	.cout());
defparam \d_writedata[29]~5 .lut_mask = 16'hAACC;
defparam \d_writedata[29]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \d_writedata[30]~6 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[30] ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[30]~6_combout ),
	.cout());
defparam \d_writedata[30]~6 .lut_mask = 16'hAACC;
defparam \d_writedata[30]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \d_writedata[31]~7 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[31] ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ),
	.datac(gnd),
	.datad(\D_ctrl_mem16~1_combout ),
	.cin(gnd),
	.combout(\d_writedata[31]~7_combout ),
	.cout());
defparam \d_writedata[31]~7 .lut_mask = 16'hAACC;
defparam \d_writedata[31]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb E_st_stall(
	.dataa(d_write1),
	.datab(\E_new_inst~q ),
	.datac(\R_ctrl_st~q ),
	.datad(av_waitrequest),
	.cin(gnd),
	.combout(\E_st_stall~combout ),
	.cout());
defparam E_st_stall.lut_mask = 16'hFFFE;
defparam E_st_stall.sum_lutc_input = "datac";

cycloneive_lcell_comb d_read_nxt(
	.dataa(d_read1),
	.datab(\E_new_inst~q ),
	.datac(\R_ctrl_ld~q ),
	.datad(WideOr11),
	.cin(gnd),
	.combout(\d_read_nxt~combout ),
	.cout());
defparam d_read_nxt.lut_mask = 16'hFFFE;
defparam d_read_nxt.sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_uncond_cti_non_br~0 (
	.dataa(\Equal0~7_combout ),
	.datab(\Equal62~11_combout ),
	.datac(\D_iw[14]~q ),
	.datad(\D_iw[15]~q ),
	.cin(gnd),
	.combout(\D_ctrl_uncond_cti_non_br~0_combout ),
	.cout());
defparam \D_ctrl_uncond_cti_non_br~0 .lut_mask = 16'hFEFF;
defparam \D_ctrl_uncond_cti_non_br~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_uncond_cti_non_br~1 (
	.dataa(\D_ctrl_jmp_direct~1_combout ),
	.datab(\D_ctrl_uncond_cti_non_br~0_combout ),
	.datac(gnd),
	.datad(\D_ctrl_force_src2_zero~3_combout ),
	.cin(gnd),
	.combout(\D_ctrl_uncond_cti_non_br~1_combout ),
	.cout());
defparam \D_ctrl_uncond_cti_non_br~1 .lut_mask = 16'hEEFF;
defparam \D_ctrl_uncond_cti_non_br~1 .sum_lutc_input = "datac";

dffeas R_ctrl_uncond_cti_non_br(
	.clk(clk_clk),
	.d(\D_ctrl_uncond_cti_non_br~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_uncond_cti_non_br~q ),
	.prn(vcc));
defparam R_ctrl_uncond_cti_non_br.is_wysiwyg = "true";
defparam R_ctrl_uncond_cti_non_br.power_up = "low";

cycloneive_lcell_comb \Equal0~19 (
	.dataa(\D_iw[5]~q ),
	.datab(\D_iw[4]~q ),
	.datac(\Equal0~5_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal0~19_combout ),
	.cout());
defparam \Equal0~19 .lut_mask = 16'hF7F7;
defparam \Equal0~19 .sum_lutc_input = "datac";

dffeas R_ctrl_br_uncond(
	.clk(clk_clk),
	.d(\Equal0~19_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_br_uncond~q ),
	.prn(vcc));
defparam R_ctrl_br_uncond.is_wysiwyg = "true";
defparam R_ctrl_br_uncond.power_up = "low";

dffeas \R_compare_op[1] (
	.clk(clk_clk),
	.d(\D_logic_op_raw[1]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_compare_op[1]~q ),
	.prn(vcc));
defparam \R_compare_op[1] .is_wysiwyg = "true";
defparam \R_compare_op[1] .power_up = "low";

cycloneive_lcell_comb \D_logic_op_raw[0]~1 (
	.dataa(\D_iw[14]~q ),
	.datab(\D_iw[3]~q ),
	.datac(\Equal0~2_combout ),
	.datad(\Equal0~3_combout ),
	.cin(gnd),
	.combout(\D_logic_op_raw[0]~1_combout ),
	.cout());
defparam \D_logic_op_raw[0]~1 .lut_mask = 16'hEFFE;
defparam \D_logic_op_raw[0]~1 .sum_lutc_input = "datac";

dffeas \R_compare_op[0] (
	.clk(clk_clk),
	.d(\D_logic_op_raw[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_compare_op[0]~q ),
	.prn(vcc));
defparam \R_compare_op[0] .is_wysiwyg = "true";
defparam \R_compare_op[0] .power_up = "low";

cycloneive_lcell_comb \Equal127~0 (
	.dataa(\E_logic_result[12]~0_combout ),
	.datab(\E_logic_result[15]~1_combout ),
	.datac(\E_logic_result[14]~2_combout ),
	.datad(\E_logic_result[13]~3_combout ),
	.cin(gnd),
	.combout(\Equal127~0_combout ),
	.cout());
defparam \Equal127~0 .lut_mask = 16'h7FFF;
defparam \Equal127~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal127~1 (
	.dataa(\E_logic_result[11]~4_combout ),
	.datab(\E_logic_result[10]~5_combout ),
	.datac(\E_logic_result[9]~6_combout ),
	.datad(\E_logic_result[8]~7_combout ),
	.cin(gnd),
	.combout(\Equal127~1_combout ),
	.cout());
defparam \Equal127~1 .lut_mask = 16'h7FFF;
defparam \Equal127~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal127~2 (
	.dataa(\E_logic_result[4]~11_combout ),
	.datab(\E_logic_result[5]~10_combout ),
	.datac(\E_logic_result[7]~8_combout ),
	.datad(\E_logic_result[6]~9_combout ),
	.cin(gnd),
	.combout(\Equal127~2_combout ),
	.cout());
defparam \Equal127~2 .lut_mask = 16'h7FFF;
defparam \Equal127~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_hi[15]~0 (
	.dataa(\D_iw[21]~q ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[31] ),
	.datac(\R_src2_use_imm~q ),
	.datad(\R_ctrl_hi_imm16~q ),
	.cin(gnd),
	.combout(\R_src2_hi[15]~0_combout ),
	.cout());
defparam \R_src2_hi[15]~0 .lut_mask = 16'hEFFE;
defparam \R_src2_hi[15]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_unsigned_lo_imm16~3 (
	.dataa(\D_iw[5]~q ),
	.datab(\Equal0~4_combout ),
	.datac(\Equal0~6_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\D_ctrl_unsigned_lo_imm16~3_combout ),
	.cout());
defparam \D_ctrl_unsigned_lo_imm16~3 .lut_mask = 16'hFAFC;
defparam \D_ctrl_unsigned_lo_imm16~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \D_ctrl_unsigned_lo_imm16~4 (
	.dataa(\D_ctrl_unsigned_lo_imm16~5_combout ),
	.datab(\D_ctrl_unsigned_lo_imm16~3_combout ),
	.datac(\D_iw[5]~q ),
	.datad(\D_ctrl_logic~0_combout ),
	.cin(gnd),
	.combout(\D_ctrl_unsigned_lo_imm16~4_combout ),
	.cout());
defparam \D_ctrl_unsigned_lo_imm16~4 .lut_mask = 16'hEFFF;
defparam \D_ctrl_unsigned_lo_imm16~4 .sum_lutc_input = "datac";

dffeas R_ctrl_unsigned_lo_imm16(
	.clk(clk_clk),
	.d(\D_ctrl_unsigned_lo_imm16~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\R_ctrl_unsigned_lo_imm16~q ),
	.prn(vcc));
defparam R_ctrl_unsigned_lo_imm16.is_wysiwyg = "true";
defparam R_ctrl_unsigned_lo_imm16.power_up = "low";

cycloneive_lcell_comb \R_src2_hi[15]~1 (
	.dataa(\R_src2_hi[15]~0_combout ),
	.datab(gnd),
	.datac(\R_ctrl_force_src2_zero~q ),
	.datad(\R_ctrl_unsigned_lo_imm16~q ),
	.cin(gnd),
	.combout(\R_src2_hi[15]~1_combout ),
	.cout());
defparam \R_src2_hi[15]~1 .lut_mask = 16'hAFFF;
defparam \R_src2_hi[15]~1 .sum_lutc_input = "datac";

dffeas \E_src2[31] (
	.clk(clk_clk),
	.d(\R_src2_hi[15]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_src2[31]~q ),
	.prn(vcc));
defparam \E_src2[31] .is_wysiwyg = "true";
defparam \E_src2[31] .power_up = "low";

cycloneive_lcell_comb \E_logic_result[31]~14 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[31]~q ),
	.datac(\E_src1[31]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[31]~14_combout ),
	.cout());
defparam \E_logic_result[31]~14 .lut_mask = 16'h6996;
defparam \E_logic_result[31]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[1]~15 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[1]~q ),
	.datac(\E_src1[1]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[1]~15_combout ),
	.cout());
defparam \E_logic_result[1]~15 .lut_mask = 16'h6996;
defparam \E_logic_result[1]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal127~3 (
	.dataa(\E_logic_result[3]~12_combout ),
	.datab(\E_logic_result[2]~13_combout ),
	.datac(\E_logic_result[31]~14_combout ),
	.datad(\E_logic_result[1]~15_combout ),
	.cin(gnd),
	.combout(\Equal127~3_combout ),
	.cout());
defparam \Equal127~3 .lut_mask = 16'h7FFF;
defparam \Equal127~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal127~4 (
	.dataa(\Equal127~0_combout ),
	.datab(\Equal127~1_combout ),
	.datac(\Equal127~2_combout ),
	.datad(\Equal127~3_combout ),
	.cin(gnd),
	.combout(\Equal127~4_combout ),
	.cout());
defparam \Equal127~4 .lut_mask = 16'hFFFE;
defparam \Equal127~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_logic_result[0]~16 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[0]~q ),
	.datac(\E_src1[0]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[0]~16_combout ),
	.cout());
defparam \E_logic_result[0]~16 .lut_mask = 16'h6996;
defparam \E_logic_result[0]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[16]~0 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[16] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[16]~0_combout ),
	.cout());
defparam \E_src2[16]~0 .lut_mask = 16'hAACC;
defparam \E_src2[16]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \R_src2_hi~2 (
	.dataa(\R_ctrl_force_src2_zero~q ),
	.datab(\R_ctrl_unsigned_lo_imm16~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\R_src2_hi~2_combout ),
	.cout());
defparam \R_src2_hi~2 .lut_mask = 16'hEEEE;
defparam \R_src2_hi~2 .sum_lutc_input = "datac";

dffeas \E_src2[16] (
	.clk(clk_clk),
	.d(\E_src2[16]~0_combout ),
	.asdata(\D_iw[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~2_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[16]~q ),
	.prn(vcc));
defparam \E_src2[16] .is_wysiwyg = "true";
defparam \E_src2[16] .power_up = "low";

cycloneive_lcell_comb \E_logic_result[16]~17 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[16]~q ),
	.datac(\E_src1[16]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[16]~17_combout ),
	.cout());
defparam \E_logic_result[16]~17 .lut_mask = 16'h6996;
defparam \E_logic_result[16]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[30]~1 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[30] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[30]~1_combout ),
	.cout());
defparam \E_src2[30]~1 .lut_mask = 16'hAACC;
defparam \E_src2[30]~1 .sum_lutc_input = "datac";

dffeas \E_src2[30] (
	.clk(clk_clk),
	.d(\E_src2[30]~1_combout ),
	.asdata(\D_iw[20]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~2_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[30]~q ),
	.prn(vcc));
defparam \E_src2[30] .is_wysiwyg = "true";
defparam \E_src2[30] .power_up = "low";

cycloneive_lcell_comb \E_logic_result[30]~18 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[30]~q ),
	.datac(\E_src1[30]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[30]~18_combout ),
	.cout());
defparam \E_logic_result[30]~18 .lut_mask = 16'h6996;
defparam \E_logic_result[30]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[29]~2 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[29] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[29]~2_combout ),
	.cout());
defparam \E_src2[29]~2 .lut_mask = 16'hAACC;
defparam \E_src2[29]~2 .sum_lutc_input = "datac";

dffeas \E_src2[29] (
	.clk(clk_clk),
	.d(\E_src2[29]~2_combout ),
	.asdata(\D_iw[19]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~2_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[29]~q ),
	.prn(vcc));
defparam \E_src2[29] .is_wysiwyg = "true";
defparam \E_src2[29] .power_up = "low";

cycloneive_lcell_comb \E_logic_result[29]~19 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[29]~q ),
	.datac(\E_src1[29]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[29]~19_combout ),
	.cout());
defparam \E_logic_result[29]~19 .lut_mask = 16'h6996;
defparam \E_logic_result[29]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal127~5 (
	.dataa(\E_logic_result[0]~16_combout ),
	.datab(\E_logic_result[16]~17_combout ),
	.datac(\E_logic_result[30]~18_combout ),
	.datad(\E_logic_result[29]~19_combout ),
	.cin(gnd),
	.combout(\Equal127~5_combout ),
	.cout());
defparam \Equal127~5 .lut_mask = 16'h7FFF;
defparam \Equal127~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[28]~3 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[28] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[28]~3_combout ),
	.cout());
defparam \E_src2[28]~3 .lut_mask = 16'hAACC;
defparam \E_src2[28]~3 .sum_lutc_input = "datac";

dffeas \E_src2[28] (
	.clk(clk_clk),
	.d(\E_src2[28]~3_combout ),
	.asdata(\D_iw[18]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~2_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[28]~q ),
	.prn(vcc));
defparam \E_src2[28] .is_wysiwyg = "true";
defparam \E_src2[28] .power_up = "low";

cycloneive_lcell_comb \E_logic_result[28]~20 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[28]~q ),
	.datac(\E_src1[28]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[28]~20_combout ),
	.cout());
defparam \E_logic_result[28]~20 .lut_mask = 16'h6996;
defparam \E_logic_result[28]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[27]~4 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[27] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[27]~4_combout ),
	.cout());
defparam \E_src2[27]~4 .lut_mask = 16'hAACC;
defparam \E_src2[27]~4 .sum_lutc_input = "datac";

dffeas \E_src2[27] (
	.clk(clk_clk),
	.d(\E_src2[27]~4_combout ),
	.asdata(\D_iw[17]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~2_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[27]~q ),
	.prn(vcc));
defparam \E_src2[27] .is_wysiwyg = "true";
defparam \E_src2[27] .power_up = "low";

cycloneive_lcell_comb \E_logic_result[27]~21 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[27]~q ),
	.datac(\E_src1[27]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[27]~21_combout ),
	.cout());
defparam \E_logic_result[27]~21 .lut_mask = 16'h6996;
defparam \E_logic_result[27]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[26]~5 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[26] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[26]~5_combout ),
	.cout());
defparam \E_src2[26]~5 .lut_mask = 16'hAACC;
defparam \E_src2[26]~5 .sum_lutc_input = "datac";

dffeas \E_src2[26] (
	.clk(clk_clk),
	.d(\E_src2[26]~5_combout ),
	.asdata(\D_iw[16]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~2_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[26]~q ),
	.prn(vcc));
defparam \E_src2[26] .is_wysiwyg = "true";
defparam \E_src2[26] .power_up = "low";

cycloneive_lcell_comb \E_logic_result[26]~22 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[26]~q ),
	.datac(\E_src1[26]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[26]~22_combout ),
	.cout());
defparam \E_logic_result[26]~22 .lut_mask = 16'h6996;
defparam \E_logic_result[26]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[25]~6 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[25] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[25]~6_combout ),
	.cout());
defparam \E_src2[25]~6 .lut_mask = 16'hAACC;
defparam \E_src2[25]~6 .sum_lutc_input = "datac";

dffeas \E_src2[25] (
	.clk(clk_clk),
	.d(\E_src2[25]~6_combout ),
	.asdata(\D_iw[15]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~2_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[25]~q ),
	.prn(vcc));
defparam \E_src2[25] .is_wysiwyg = "true";
defparam \E_src2[25] .power_up = "low";

cycloneive_lcell_comb \E_logic_result[25]~23 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[25]~q ),
	.datac(\E_src1[25]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[25]~23_combout ),
	.cout());
defparam \E_logic_result[25]~23 .lut_mask = 16'h6996;
defparam \E_logic_result[25]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal127~6 (
	.dataa(\E_logic_result[28]~20_combout ),
	.datab(\E_logic_result[27]~21_combout ),
	.datac(\E_logic_result[26]~22_combout ),
	.datad(\E_logic_result[25]~23_combout ),
	.cin(gnd),
	.combout(\Equal127~6_combout ),
	.cout());
defparam \Equal127~6 .lut_mask = 16'h7FFF;
defparam \Equal127~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[24]~7 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[24] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[24]~7_combout ),
	.cout());
defparam \E_src2[24]~7 .lut_mask = 16'hAACC;
defparam \E_src2[24]~7 .sum_lutc_input = "datac";

dffeas \E_src2[24] (
	.clk(clk_clk),
	.d(\E_src2[24]~7_combout ),
	.asdata(\D_iw[14]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~2_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[24]~q ),
	.prn(vcc));
defparam \E_src2[24] .is_wysiwyg = "true";
defparam \E_src2[24] .power_up = "low";

cycloneive_lcell_comb \E_logic_result[24]~24 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[24]~q ),
	.datac(\E_src1[24]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[24]~24_combout ),
	.cout());
defparam \E_logic_result[24]~24 .lut_mask = 16'h6996;
defparam \E_logic_result[24]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[23]~8 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[23] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[23]~8_combout ),
	.cout());
defparam \E_src2[23]~8 .lut_mask = 16'hAACC;
defparam \E_src2[23]~8 .sum_lutc_input = "datac";

dffeas \E_src2[23] (
	.clk(clk_clk),
	.d(\E_src2[23]~8_combout ),
	.asdata(\D_iw[13]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~2_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[23]~q ),
	.prn(vcc));
defparam \E_src2[23] .is_wysiwyg = "true";
defparam \E_src2[23] .power_up = "low";

cycloneive_lcell_comb \E_logic_result[23]~25 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[23]~q ),
	.datac(\E_src1[23]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[23]~25_combout ),
	.cout());
defparam \E_logic_result[23]~25 .lut_mask = 16'h6996;
defparam \E_logic_result[23]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[22]~9 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[22] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[22]~9_combout ),
	.cout());
defparam \E_src2[22]~9 .lut_mask = 16'hAACC;
defparam \E_src2[22]~9 .sum_lutc_input = "datac";

dffeas \E_src2[22] (
	.clk(clk_clk),
	.d(\E_src2[22]~9_combout ),
	.asdata(\D_iw[12]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~2_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[22]~q ),
	.prn(vcc));
defparam \E_src2[22] .is_wysiwyg = "true";
defparam \E_src2[22] .power_up = "low";

cycloneive_lcell_comb \E_logic_result[22]~26 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[22]~q ),
	.datac(\E_src1[22]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[22]~26_combout ),
	.cout());
defparam \E_logic_result[22]~26 .lut_mask = 16'h6996;
defparam \E_logic_result[22]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[21]~10 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[21] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[21]~10_combout ),
	.cout());
defparam \E_src2[21]~10 .lut_mask = 16'hAACC;
defparam \E_src2[21]~10 .sum_lutc_input = "datac";

dffeas \E_src2[21] (
	.clk(clk_clk),
	.d(\E_src2[21]~10_combout ),
	.asdata(\D_iw[11]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~2_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[21]~q ),
	.prn(vcc));
defparam \E_src2[21] .is_wysiwyg = "true";
defparam \E_src2[21] .power_up = "low";

cycloneive_lcell_comb \E_logic_result[21]~27 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[21]~q ),
	.datac(\E_src1[21]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[21]~27_combout ),
	.cout());
defparam \E_logic_result[21]~27 .lut_mask = 16'h6996;
defparam \E_logic_result[21]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal127~7 (
	.dataa(\E_logic_result[24]~24_combout ),
	.datab(\E_logic_result[23]~25_combout ),
	.datac(\E_logic_result[22]~26_combout ),
	.datad(\E_logic_result[21]~27_combout ),
	.cin(gnd),
	.combout(\Equal127~7_combout ),
	.cout());
defparam \Equal127~7 .lut_mask = 16'h7FFF;
defparam \Equal127~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[20]~11 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[20] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[20]~11_combout ),
	.cout());
defparam \E_src2[20]~11 .lut_mask = 16'hAACC;
defparam \E_src2[20]~11 .sum_lutc_input = "datac";

dffeas \E_src2[20] (
	.clk(clk_clk),
	.d(\E_src2[20]~11_combout ),
	.asdata(\D_iw[10]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~2_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[20]~q ),
	.prn(vcc));
defparam \E_src2[20] .is_wysiwyg = "true";
defparam \E_src2[20] .power_up = "low";

cycloneive_lcell_comb \E_logic_result[20]~28 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[20]~q ),
	.datac(\E_src1[20]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[20]~28_combout ),
	.cout());
defparam \E_logic_result[20]~28 .lut_mask = 16'h6996;
defparam \E_logic_result[20]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[19]~12 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[19] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[19]~12_combout ),
	.cout());
defparam \E_src2[19]~12 .lut_mask = 16'hAACC;
defparam \E_src2[19]~12 .sum_lutc_input = "datac";

dffeas \E_src2[19] (
	.clk(clk_clk),
	.d(\E_src2[19]~12_combout ),
	.asdata(\D_iw[9]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~2_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[19]~q ),
	.prn(vcc));
defparam \E_src2[19] .is_wysiwyg = "true";
defparam \E_src2[19] .power_up = "low";

cycloneive_lcell_comb \E_logic_result[19]~29 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[19]~q ),
	.datac(\E_src1[19]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[19]~29_combout ),
	.cout());
defparam \E_logic_result[19]~29 .lut_mask = 16'h6996;
defparam \E_logic_result[19]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[18]~13 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[18] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[18]~13_combout ),
	.cout());
defparam \E_src2[18]~13 .lut_mask = 16'hAACC;
defparam \E_src2[18]~13 .sum_lutc_input = "datac";

dffeas \E_src2[18] (
	.clk(clk_clk),
	.d(\E_src2[18]~13_combout ),
	.asdata(\D_iw[8]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~2_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[18]~q ),
	.prn(vcc));
defparam \E_src2[18] .is_wysiwyg = "true";
defparam \E_src2[18] .power_up = "low";

cycloneive_lcell_comb \E_logic_result[18]~30 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[18]~q ),
	.datac(\E_src1[18]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[18]~30_combout ),
	.cout());
defparam \E_logic_result[18]~30 .lut_mask = 16'h6996;
defparam \E_logic_result[18]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_src2[17]~14 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[17] ),
	.datab(\D_iw[21]~q ),
	.datac(gnd),
	.datad(\R_src2_use_imm~q ),
	.cin(gnd),
	.combout(\E_src2[17]~14_combout ),
	.cout());
defparam \E_src2[17]~14 .lut_mask = 16'hAACC;
defparam \E_src2[17]~14 .sum_lutc_input = "datac";

dffeas \E_src2[17] (
	.clk(clk_clk),
	.d(\E_src2[17]~14_combout ),
	.asdata(\D_iw[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\R_src2_hi~2_combout ),
	.sload(\R_ctrl_hi_imm16~q ),
	.ena(vcc),
	.q(\E_src2[17]~q ),
	.prn(vcc));
defparam \E_src2[17] .is_wysiwyg = "true";
defparam \E_src2[17] .power_up = "low";

cycloneive_lcell_comb \E_logic_result[17]~31 (
	.dataa(\R_logic_op[1]~q ),
	.datab(\E_src2[17]~q ),
	.datac(\E_src1[17]~q ),
	.datad(\R_logic_op[0]~q ),
	.cin(gnd),
	.combout(\E_logic_result[17]~31_combout ),
	.cout());
defparam \E_logic_result[17]~31 .lut_mask = 16'h6996;
defparam \E_logic_result[17]~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal127~8 (
	.dataa(\E_logic_result[20]~28_combout ),
	.datab(\E_logic_result[19]~29_combout ),
	.datac(\E_logic_result[18]~30_combout ),
	.datad(\E_logic_result[17]~31_combout ),
	.cin(gnd),
	.combout(\Equal127~8_combout ),
	.cout());
defparam \Equal127~8 .lut_mask = 16'h7FFF;
defparam \Equal127~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal127~9 (
	.dataa(\Equal127~5_combout ),
	.datab(\Equal127~6_combout ),
	.datac(\Equal127~7_combout ),
	.datad(\Equal127~8_combout ),
	.cin(gnd),
	.combout(\Equal127~9_combout ),
	.cout());
defparam \Equal127~9 .lut_mask = 16'hFFFE;
defparam \Equal127~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_cmp_result~0 (
	.dataa(\R_compare_op[1]~q ),
	.datab(\R_compare_op[0]~q ),
	.datac(\Equal127~4_combout ),
	.datad(\Equal127~9_combout ),
	.cin(gnd),
	.combout(\E_cmp_result~0_combout ),
	.cout());
defparam \E_cmp_result~0 .lut_mask = 16'h6996;
defparam \E_cmp_result~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_invert_arith_src_msb~1 (
	.dataa(\Equal0~7_combout ),
	.datab(\Equal62~0_combout ),
	.datac(\D_iw[15]~q ),
	.datad(\D_iw[14]~q ),
	.cin(gnd),
	.combout(\E_invert_arith_src_msb~1_combout ),
	.cout());
defparam \E_invert_arith_src_msb~1 .lut_mask = 16'hEFFE;
defparam \E_invert_arith_src_msb~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_invert_arith_src_msb~2 (
	.dataa(\R_valid~q ),
	.datab(\E_invert_arith_src_msb~1_combout ),
	.datac(\D_iw[5]~q ),
	.datad(\E_invert_arith_src_msb~0_combout ),
	.cin(gnd),
	.combout(\E_invert_arith_src_msb~2_combout ),
	.cout());
defparam \E_invert_arith_src_msb~2 .lut_mask = 16'hEFFF;
defparam \E_invert_arith_src_msb~2 .sum_lutc_input = "datac";

dffeas E_invert_arith_src_msb(
	.clk(clk_clk),
	.d(\E_invert_arith_src_msb~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\E_invert_arith_src_msb~q ),
	.prn(vcc));
defparam E_invert_arith_src_msb.is_wysiwyg = "true";
defparam E_invert_arith_src_msb.power_up = "low";

cycloneive_lcell_comb \Add1~50 (
	.dataa(\E_alu_sub~q ),
	.datab(\E_src2[31]~q ),
	.datac(\E_invert_arith_src_msb~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Add1~50_combout ),
	.cout());
defparam \Add1~50 .lut_mask = 16'h9696;
defparam \Add1~50 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_arith_src1[31] (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_invert_arith_src_msb~q ),
	.datad(\E_src1[31]~q ),
	.cin(gnd),
	.combout(\E_arith_src1[31]~combout ),
	.cout());
defparam \E_arith_src1[31] .lut_mask = 16'h0FF0;
defparam \E_arith_src1[31] .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~51 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[30]~q ),
	.cin(gnd),
	.combout(\Add1~51_combout ),
	.cout());
defparam \Add1~51 .lut_mask = 16'h0FF0;
defparam \Add1~51 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~52 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[29]~q ),
	.cin(gnd),
	.combout(\Add1~52_combout ),
	.cout());
defparam \Add1~52 .lut_mask = 16'h0FF0;
defparam \Add1~52 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[28]~q ),
	.cin(gnd),
	.combout(\Add1~53_combout ),
	.cout());
defparam \Add1~53 .lut_mask = 16'h0FF0;
defparam \Add1~53 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~54 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[27]~q ),
	.cin(gnd),
	.combout(\Add1~54_combout ),
	.cout());
defparam \Add1~54 .lut_mask = 16'h0FF0;
defparam \Add1~54 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~55 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[26]~q ),
	.cin(gnd),
	.combout(\Add1~55_combout ),
	.cout());
defparam \Add1~55 .lut_mask = 16'h0FF0;
defparam \Add1~55 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~56 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[25]~q ),
	.cin(gnd),
	.combout(\Add1~56_combout ),
	.cout());
defparam \Add1~56 .lut_mask = 16'h0FF0;
defparam \Add1~56 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[24]~q ),
	.cin(gnd),
	.combout(\Add1~57_combout ),
	.cout());
defparam \Add1~57 .lut_mask = 16'h0FF0;
defparam \Add1~57 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~58 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[23]~q ),
	.cin(gnd),
	.combout(\Add1~58_combout ),
	.cout());
defparam \Add1~58 .lut_mask = 16'h0FF0;
defparam \Add1~58 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~59 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[22]~q ),
	.cin(gnd),
	.combout(\Add1~59_combout ),
	.cout());
defparam \Add1~59 .lut_mask = 16'h0FF0;
defparam \Add1~59 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~60 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[21]~q ),
	.cin(gnd),
	.combout(\Add1~60_combout ),
	.cout());
defparam \Add1~60 .lut_mask = 16'h0FF0;
defparam \Add1~60 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[20]~q ),
	.cin(gnd),
	.combout(\Add1~61_combout ),
	.cout());
defparam \Add1~61 .lut_mask = 16'h0FF0;
defparam \Add1~61 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~62 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[19]~q ),
	.cin(gnd),
	.combout(\Add1~62_combout ),
	.cout());
defparam \Add1~62 .lut_mask = 16'h0FF0;
defparam \Add1~62 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~63 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[18]~q ),
	.cin(gnd),
	.combout(\Add1~63_combout ),
	.cout());
defparam \Add1~63 .lut_mask = 16'h0FF0;
defparam \Add1~63 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~64 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[17]~q ),
	.cin(gnd),
	.combout(\Add1~64_combout ),
	.cout());
defparam \Add1~64 .lut_mask = 16'h0FF0;
defparam \Add1~64 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\E_alu_sub~q ),
	.datad(\E_src2[16]~q ),
	.cin(gnd),
	.combout(\Add1~65_combout ),
	.cout());
defparam \Add1~65 .lut_mask = 16'h0FF0;
defparam \Add1~65 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~98 (
	.dataa(\E_alu_sub~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add1~97 ),
	.combout(\Add1~98_combout ),
	.cout());
defparam \Add1~98 .lut_mask = 16'h5A5A;
defparam \Add1~98 .sum_lutc_input = "cin";

cycloneive_lcell_comb \E_cmp_result~1 (
	.dataa(\E_cmp_result~0_combout ),
	.datab(\R_compare_op[1]~q ),
	.datac(\Add1~98_combout ),
	.datad(\R_compare_op[0]~q ),
	.cin(gnd),
	.combout(\E_cmp_result~1_combout ),
	.cout());
defparam \E_cmp_result~1 .lut_mask = 16'hEBBE;
defparam \E_cmp_result~1 .sum_lutc_input = "datac";

dffeas W_cmp_result(
	.clk(clk_clk),
	.d(\E_cmp_result~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_cmp_result~q ),
	.prn(vcc));
defparam W_cmp_result.is_wysiwyg = "true";
defparam W_cmp_result.power_up = "low";

cycloneive_lcell_comb \F_pc_sel_nxt~0 (
	.dataa(\R_ctrl_uncond_cti_non_br~q ),
	.datab(\R_ctrl_br_uncond~q ),
	.datac(\W_cmp_result~q ),
	.datad(\R_ctrl_br~q ),
	.cin(gnd),
	.combout(\F_pc_sel_nxt~0_combout ),
	.cout());
defparam \F_pc_sel_nxt~0 .lut_mask = 16'hFFFE;
defparam \F_pc_sel_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[10]~0 (
	.dataa(\Add1~39_combout ),
	.datab(\F_pc_plus_one[10]~20_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[10]~0_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[10]~0 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[10]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[9]~1 (
	.dataa(\F_pc_sel_nxt~0_combout ),
	.datab(\F_pc_sel_nxt.10~0_combout ),
	.datac(\F_pc_plus_one[9]~18_combout ),
	.datad(\Add1~37_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[9]~1_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[9]~1 .lut_mask = 16'hFFF6;
defparam \F_pc_no_crst_nxt[9]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[9]~2 (
	.dataa(\R_ctrl_break~q ),
	.datab(\R_ctrl_exception~q ),
	.datac(\F_pc_no_crst_nxt[9]~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[9]~2_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[9]~2 .lut_mask = 16'hFBFB;
defparam \F_pc_no_crst_nxt[9]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[8]~3 (
	.dataa(\Add1~35_combout ),
	.datab(\F_pc_plus_one[8]~16_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[8]~3_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[8]~3 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[8]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[7]~4 (
	.dataa(\Add1~33_combout ),
	.datab(\F_pc_plus_one[7]~14_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[7]~4_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[7]~4 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[7]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[6]~5 (
	.dataa(\Add1~31_combout ),
	.datab(\F_pc_plus_one[6]~12_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[6]~5_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[6]~5 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[6]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[5]~6 (
	.dataa(\Add1~29_combout ),
	.datab(\F_pc_plus_one[5]~10_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[5]~6_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[5]~6 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[5]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[4]~7 (
	.dataa(\Add1~27_combout ),
	.datab(\F_pc_plus_one[4]~8_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[4]~7_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[4]~7 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[4]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[3]~8 (
	.dataa(\F_pc_sel_nxt.10~0_combout ),
	.datab(\Add1~25_combout ),
	.datac(\F_pc_plus_one[3]~6_combout ),
	.datad(\F_pc_sel_nxt~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[3]~8_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[3]~8 .lut_mask = 16'hFAFC;
defparam \F_pc_no_crst_nxt[3]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[2]~9 (
	.dataa(\Add1~23_combout ),
	.datab(\F_pc_plus_one[2]~4_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[2]~9_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[2]~9 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[2]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[1]~10 (
	.dataa(\Add1~21_combout ),
	.datab(\F_pc_plus_one[1]~2_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[1]~10_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[1]~10 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[1]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[0]~11 (
	.dataa(\Add1~19_combout ),
	.datab(\F_pc_plus_one[0]~0_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[0]~11_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[0]~11 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[0]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[13]~12 (
	.dataa(\R_ctrl_break~q ),
	.datab(\F_pc_plus_one[13]~26_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\R_ctrl_exception~q ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[13]~12_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[13]~12 .lut_mask = 16'hEFFF;
defparam \F_pc_no_crst_nxt[13]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[13]~13 (
	.dataa(\F_pc_no_crst_nxt[13]~12_combout ),
	.datab(\Add1~48_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\R_ctrl_exception~q ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[13]~13_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[13]~13 .lut_mask = 16'hFEFF;
defparam \F_pc_no_crst_nxt[13]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[12]~14 (
	.dataa(\Add1~46_combout ),
	.datab(\F_pc_plus_one[12]~24_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[12]~14_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[12]~14 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[12]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \F_pc_no_crst_nxt[11]~15 (
	.dataa(\Add1~44_combout ),
	.datab(\F_pc_plus_one[11]~22_combout ),
	.datac(\F_pc_sel_nxt~0_combout ),
	.datad(\F_pc_sel_nxt.10~0_combout ),
	.cin(gnd),
	.combout(\F_pc_no_crst_nxt[11]~15_combout ),
	.cout());
defparam \F_pc_no_crst_nxt[11]~15 .lut_mask = 16'hACFF;
defparam \F_pc_no_crst_nxt[11]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \i_read_nxt~0 (
	.dataa(\W_valid~q ),
	.datab(i_read1),
	.datac(src1_valid),
	.datad(read_latency_shift_reg_05),
	.cin(gnd),
	.combout(\i_read_nxt~0_combout ),
	.cout());
defparam \i_read_nxt~0 .lut_mask = 16'hFFFD;
defparam \i_read_nxt~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \hbreak_enabled~0 (
	.dataa(\D_op_cmpge~0_combout ),
	.datab(\Equal62~9_combout ),
	.datac(hbreak_enabled1),
	.datad(\R_ctrl_break~q ),
	.cin(gnd),
	.combout(\hbreak_enabled~0_combout ),
	.cout());
defparam \hbreak_enabled~0 .lut_mask = 16'hFFF7;
defparam \hbreak_enabled~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_mem_byte_en[0]~0 (
	.dataa(\D_ctrl_mem16~1_combout ),
	.datab(\D_ctrl_mem8~1_combout ),
	.datac(\Add1~15_combout ),
	.datad(\Add1~17_combout ),
	.cin(gnd),
	.combout(\E_mem_byte_en[0]~0_combout ),
	.cout());
defparam \E_mem_byte_en[0]~0 .lut_mask = 16'h6FFF;
defparam \E_mem_byte_en[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \d_byteenable[3]~0 (
	.dataa(\D_ctrl_mem16~0_combout ),
	.datab(\D_ctrl_mem8~0_combout ),
	.datac(gnd),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\d_byteenable[3]~0_combout ),
	.cout());
defparam \d_byteenable[3]~0 .lut_mask = 16'hEEFF;
defparam \d_byteenable[3]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[22]~0 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[22] ),
	.datac(gnd),
	.datad(\d_byteenable[3]~0_combout ),
	.cin(gnd),
	.combout(\E_st_data[22]~0_combout ),
	.cout());
defparam \E_st_data[22]~0 .lut_mask = 16'hAACC;
defparam \E_st_data[22]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_mem_byte_en[2]~1 (
	.dataa(\D_ctrl_mem16~1_combout ),
	.datab(\Add1~17_combout ),
	.datac(\D_ctrl_mem8~1_combout ),
	.datad(\Add1~15_combout ),
	.cin(gnd),
	.combout(\E_mem_byte_en[2]~1_combout ),
	.cout());
defparam \E_mem_byte_en[2]~1 .lut_mask = 16'hDEFF;
defparam \E_mem_byte_en[2]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[23]~1 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[23] ),
	.datac(gnd),
	.datad(\d_byteenable[3]~0_combout ),
	.cin(gnd),
	.combout(\E_st_data[23]~1_combout ),
	.cout());
defparam \E_st_data[23]~1 .lut_mask = 16'hAACC;
defparam \E_st_data[23]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_mem_byte_en[3]~2 (
	.dataa(\D_ctrl_mem16~1_combout ),
	.datab(\Add1~17_combout ),
	.datac(\Add1~15_combout ),
	.datad(\D_ctrl_mem8~1_combout ),
	.cin(gnd),
	.combout(\E_mem_byte_en[3]~2_combout ),
	.cout());
defparam \E_mem_byte_en[3]~2 .lut_mask = 16'hFDFE;
defparam \E_mem_byte_en[3]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[11]~2 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[11]~2_combout ),
	.cout());
defparam \E_st_data[11]~2 .lut_mask = 16'hEFFE;
defparam \E_st_data[11]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_mem_byte_en[1]~3 (
	.dataa(\D_ctrl_mem16~1_combout ),
	.datab(\D_ctrl_mem8~1_combout ),
	.datac(\Add1~15_combout ),
	.datad(\Add1~17_combout ),
	.cin(gnd),
	.combout(\E_mem_byte_en[1]~3_combout ),
	.cout());
defparam \E_mem_byte_en[1]~3 .lut_mask = 16'hF6FF;
defparam \E_mem_byte_en[1]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[13]~3 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[13]~3_combout ),
	.cout());
defparam \E_st_data[13]~3 .lut_mask = 16'hEFFE;
defparam \E_st_data[13]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[16]~4 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[16] ),
	.datac(gnd),
	.datad(\d_byteenable[3]~0_combout ),
	.cin(gnd),
	.combout(\E_st_data[16]~4_combout ),
	.cout());
defparam \E_st_data[16]~4 .lut_mask = 16'hAACC;
defparam \E_st_data[16]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[12]~5 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[12]~5_combout ),
	.cout());
defparam \E_st_data[12]~5 .lut_mask = 16'hEFFE;
defparam \E_st_data[12]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[14]~6 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[14]~6_combout ),
	.cout());
defparam \E_st_data[14]~6 .lut_mask = 16'hEFFE;
defparam \E_st_data[14]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[15]~7 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[15]~7_combout ),
	.cout());
defparam \E_st_data[15]~7 .lut_mask = 16'hEFFE;
defparam \E_st_data[15]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[18]~8 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[18] ),
	.datac(gnd),
	.datad(\d_byteenable[3]~0_combout ),
	.cin(gnd),
	.combout(\E_st_data[18]~8_combout ),
	.cout());
defparam \E_st_data[18]~8 .lut_mask = 16'hAACC;
defparam \E_st_data[18]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[17]~9 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[17] ),
	.datac(gnd),
	.datad(\d_byteenable[3]~0_combout ),
	.cin(gnd),
	.combout(\E_st_data[17]~9_combout ),
	.cout());
defparam \E_st_data[17]~9 .lut_mask = 16'hAACC;
defparam \E_st_data[17]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[10]~10 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[10]~10_combout ),
	.cout());
defparam \E_st_data[10]~10 .lut_mask = 16'hEFFE;
defparam \E_st_data[10]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[9]~11 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[9]~11_combout ),
	.cout());
defparam \E_st_data[9]~11 .lut_mask = 16'hEFFE;
defparam \E_st_data[9]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[8]~12 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.datac(\D_ctrl_mem8~0_combout ),
	.datad(\D_iw[4]~q ),
	.cin(gnd),
	.combout(\E_st_data[8]~12_combout ),
	.cout());
defparam \E_st_data[8]~12 .lut_mask = 16'hEFFE;
defparam \E_st_data[8]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[21]~13 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[21] ),
	.datac(gnd),
	.datad(\d_byteenable[3]~0_combout ),
	.cin(gnd),
	.combout(\E_st_data[21]~13_combout ),
	.cout());
defparam \E_st_data[21]~13 .lut_mask = 16'hAACC;
defparam \E_st_data[21]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[19]~14 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[19] ),
	.datac(gnd),
	.datad(\d_byteenable[3]~0_combout ),
	.cin(gnd),
	.combout(\E_st_data[19]~14_combout ),
	.cout());
defparam \E_st_data[19]~14 .lut_mask = 16'hAACC;
defparam \E_st_data[19]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \E_st_data[20]~15 (
	.dataa(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.datab(\nios_mcu_nios_cpu_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[20] ),
	.datac(gnd),
	.datad(\d_byteenable[3]~0_combout ),
	.cin(gnd),
	.combout(\E_st_data[20]~15_combout ),
	.cout());
defparam \E_st_data[20]~15 .lut_mask = 16'hAACC;
defparam \E_st_data[20]~15 .sum_lutc_input = "datac";

endmodule

module nios_mcu_nios_mcu_nios_cpu_cpu_nios2_oci (
	sr_0,
	jtag_break,
	readdata_0,
	readdata_1,
	readdata_3,
	readdata_2,
	ir_out_0,
	ir_out_1,
	r_sync_rst,
	m0_write,
	saved_grant_0,
	waitrequest,
	mem_used_1,
	WideOr1,
	rf_source_valid,
	hbreak_enabled,
	address_nxt,
	r_early_rst,
	oci_ienable_0,
	oci_single_step_mode,
	readdata_22,
	readdata_23,
	readdata_24,
	readdata_25,
	readdata_26,
	readdata_11,
	readdata_13,
	readdata_16,
	readdata_12,
	readdata_5,
	readdata_4,
	readdata_14,
	readdata_15,
	readdata_18,
	readdata_17,
	readdata_10,
	readdata_9,
	readdata_8,
	readdata_7,
	readdata_6,
	readdata_21,
	readdata_19,
	readdata_20,
	debugaccess_nxt,
	writedata_nxt,
	byteenable_nxt,
	readdata_27,
	readdata_28,
	readdata_29,
	readdata_30,
	readdata_31,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	sr_0;
output 	jtag_break;
output 	readdata_0;
output 	readdata_1;
output 	readdata_3;
output 	readdata_2;
output 	ir_out_0;
output 	ir_out_1;
input 	r_sync_rst;
input 	m0_write;
input 	saved_grant_0;
output 	waitrequest;
input 	mem_used_1;
input 	WideOr1;
input 	rf_source_valid;
input 	hbreak_enabled;
input 	[8:0] address_nxt;
input 	r_early_rst;
output 	oci_ienable_0;
output 	oci_single_step_mode;
output 	readdata_22;
output 	readdata_23;
output 	readdata_24;
output 	readdata_25;
output 	readdata_26;
output 	readdata_11;
output 	readdata_13;
output 	readdata_16;
output 	readdata_12;
output 	readdata_5;
output 	readdata_4;
output 	readdata_14;
output 	readdata_15;
output 	readdata_18;
output 	readdata_17;
output 	readdata_10;
output 	readdata_9;
output 	readdata_8;
output 	readdata_7;
output 	readdata_6;
output 	readdata_21;
output 	readdata_19;
output 	readdata_20;
input 	debugaccess_nxt;
input 	[31:0] writedata_nxt;
input 	[3:0] byteenable_nxt;
output 	readdata_27;
output 	readdata_28;
output 	readdata_29;
output 	readdata_30;
output 	readdata_31;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[0] ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[1] ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[2] ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[22] ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[23] ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[24] ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[25] ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[26] ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[11] ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[13] ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[16] ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[12] ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[3] ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[5] ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[4] ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[14] ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[15] ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[18] ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[17] ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[10] ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[9] ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[8] ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[7] ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[6] ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[21] ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[19] ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[20] ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[4]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[12]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[5]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[18]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[27] ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[28] ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[29] ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[30] ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[31] ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[8]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[29]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[0]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[0]~q ;
wire \write~q ;
wire \read~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[1]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[1]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[0]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[36]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[37]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|ir[0]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|ir[1]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|enable_action_strobe~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[3]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[35]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|take_action_ocimem_b~combout ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~0_combout ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci_debug|monitor_ready~q ;
wire \write~0_combout ;
wire \write~1_combout ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[17]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~1_combout ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[34]~q ;
wire \read~0_combout ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[2]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[2]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[1]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[4]~q ;
wire \debugaccess~q ;
wire \writedata[0]~q ;
wire \address[0]~q ;
wire \address[1]~q ;
wire \address[2]~q ;
wire \address[3]~q ;
wire \address[4]~q ;
wire \address[5]~q ;
wire \address[6]~q ;
wire \address[7]~q ;
wire \byteenable[0]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|Equal0~2_combout ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|take_action_ocireg~0_combout ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[25]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[21]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[20]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~combout ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[33]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[32]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[31]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[30]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[29]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[28]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[27]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[26]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[3]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[3]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[2]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[5]~q ;
wire \writedata[1]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci_debug|monitor_error~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|Equal1~0_combout ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_reg_readdata[0]~0_combout ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[19]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[18]~q ;
wire \writedata[3]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_ienable[16]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci_debug|monitor_go~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[16]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[16]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[4]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[6]~q ;
wire \writedata[2]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[24]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[24]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[20]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[20]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[19]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[19]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[22]~q ;
wire \writedata[22]~q ;
wire \byteenable[2]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[23]~q ;
wire \writedata[23]~q ;
wire \writedata[24]~q ;
wire \byteenable[3]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[25]~q ;
wire \writedata[25]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[26]~q ;
wire \writedata[26]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[11]~q ;
wire \writedata[11]~q ;
wire \byteenable[1]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[13]~q ;
wire \writedata[13]~q ;
wire \writedata[16]~q ;
wire \writedata[12]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[23]~q ;
wire \writedata[5]~q ;
wire \writedata[4]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[14]~q ;
wire \writedata[14]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[15]~q ;
wire \writedata[15]~q ;
wire \writedata[18]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[17]~q ;
wire \writedata[17]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[10]~q ;
wire \writedata[10]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[9]~q ;
wire \writedata[9]~q ;
wire \writedata[8]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[7]~q ;
wire \writedata[7]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[6]~q ;
wire \writedata[6]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[21]~q ;
wire \writedata[21]~q ;
wire \writedata[19]~q ;
wire \writedata[20]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[17]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[16]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci_debug|resetlatch~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[31]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[31]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[30]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[30]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[29]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[28]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[28]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[27]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[27]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[26]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[25]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[5]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[7]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[24]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[18]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[21]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[22]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[14]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[15]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[8]~q ;
wire \writedata[27]~q ;
wire \writedata[28]~q ;
wire \writedata[29]~q ;
wire \writedata[30]~q ;
wire \writedata[31]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[13]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[12]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[11]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[10]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[9]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[6]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[22]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[15]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[7]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[23]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[13]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[14]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[12]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[11]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[10]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[9]~q ;
wire \the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[8]~q ;
wire \address[8]~q ;
wire \readdata~9_combout ;
wire \readdata~10_combout ;
wire \readdata~11_combout ;
wire \readdata~0_combout ;
wire \readdata~1_combout ;
wire \readdata~2_combout ;
wire \readdata~3_combout ;
wire \readdata~4_combout ;
wire \readdata~5_combout ;
wire \readdata~6_combout ;
wire \readdata~7_combout ;
wire \readdata~8_combout ;
wire \readdata~12_combout ;
wire \readdata~13_combout ;
wire \readdata~14_combout ;
wire \readdata~15_combout ;
wire \readdata~16_combout ;
wire \readdata~17_combout ;
wire \readdata~18_combout ;
wire \readdata~19_combout ;
wire \readdata~20_combout ;
wire \readdata~21_combout ;
wire \readdata~22_combout ;
wire \readdata~23_combout ;
wire \readdata~24_combout ;
wire \readdata~25_combout ;
wire \readdata~26_combout ;
wire \readdata~27_combout ;
wire \readdata~28_combout ;
wire \readdata~29_combout ;
wire \readdata~30_combout ;


nios_mcu_nios_mcu_nios_cpu_cpu_debug_slave_wrapper the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper(
	.sr_0(sr_0),
	.MonDReg_4(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[4]~q ),
	.MonDReg_12(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[12]~q ),
	.MonDReg_5(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[5]~q ),
	.MonDReg_18(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[18]~q ),
	.MonDReg_8(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[8]~q ),
	.MonDReg_29(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[29]~q ),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.break_readreg_0(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[0]~q ),
	.MonDReg_0(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[0]~q ),
	.break_readreg_1(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[1]~q ),
	.MonDReg_1(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[1]~q ),
	.jdo_0(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[0]~q ),
	.jdo_36(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[36]~q ),
	.jdo_37(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[37]~q ),
	.ir_0(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|ir[0]~q ),
	.ir_1(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|ir[1]~q ),
	.enable_action_strobe(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|enable_action_strobe~q ),
	.jdo_3(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[3]~q ),
	.jdo_35(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[35]~q ),
	.take_action_ocimem_b(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|take_action_ocimem_b~combout ),
	.take_action_ocimem_a(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~0_combout ),
	.monitor_ready(\the_nios_mcu_nios_cpu_cpu_nios2_oci_debug|monitor_ready~q ),
	.hbreak_enabled(hbreak_enabled),
	.jdo_17(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[17]~q ),
	.take_action_ocimem_a1(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~1_combout ),
	.jdo_34(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[34]~q ),
	.break_readreg_2(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[2]~q ),
	.MonDReg_2(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[2]~q ),
	.jdo_1(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[1]~q ),
	.jdo_4(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[4]~q ),
	.jdo_25(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[25]~q ),
	.jdo_21(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[21]~q ),
	.jdo_20(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[20]~q ),
	.take_action_ocimem_a2(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~combout ),
	.jdo_33(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[33]~q ),
	.jdo_32(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[32]~q ),
	.jdo_31(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[31]~q ),
	.jdo_30(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[30]~q ),
	.jdo_29(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[29]~q ),
	.jdo_28(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[28]~q ),
	.jdo_27(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[27]~q ),
	.jdo_26(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[26]~q ),
	.break_readreg_3(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[3]~q ),
	.MonDReg_3(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[3]~q ),
	.jdo_2(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[2]~q ),
	.jdo_5(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[5]~q ),
	.monitor_error(\the_nios_mcu_nios_cpu_cpu_nios2_oci_debug|monitor_error~q ),
	.jdo_19(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[19]~q ),
	.jdo_18(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[18]~q ),
	.break_readreg_16(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[16]~q ),
	.MonDReg_16(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[16]~q ),
	.break_readreg_4(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[4]~q ),
	.jdo_6(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[6]~q ),
	.break_readreg_24(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[24]~q ),
	.MonDReg_24(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[24]~q ),
	.break_readreg_20(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[20]~q ),
	.MonDReg_20(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[20]~q ),
	.break_readreg_19(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[19]~q ),
	.MonDReg_19(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[19]~q ),
	.MonDReg_22(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[22]~q ),
	.MonDReg_23(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[23]~q ),
	.MonDReg_25(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[25]~q ),
	.MonDReg_26(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[26]~q ),
	.MonDReg_11(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[11]~q ),
	.MonDReg_13(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[13]~q ),
	.jdo_23(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[23]~q ),
	.MonDReg_14(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[14]~q ),
	.MonDReg_15(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[15]~q ),
	.MonDReg_17(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[17]~q ),
	.MonDReg_10(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[10]~q ),
	.MonDReg_9(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[9]~q ),
	.MonDReg_7(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[7]~q ),
	.MonDReg_6(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[6]~q ),
	.MonDReg_21(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[21]~q ),
	.break_readreg_17(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[17]~q ),
	.jdo_16(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[16]~q ),
	.resetlatch(\the_nios_mcu_nios_cpu_cpu_nios2_oci_debug|resetlatch~q ),
	.break_readreg_31(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[31]~q ),
	.MonDReg_31(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[31]~q ),
	.break_readreg_30(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[30]~q ),
	.MonDReg_30(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[30]~q ),
	.break_readreg_29(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[29]~q ),
	.break_readreg_28(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[28]~q ),
	.MonDReg_28(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[28]~q ),
	.break_readreg_27(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[27]~q ),
	.MonDReg_27(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[27]~q ),
	.break_readreg_26(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[26]~q ),
	.break_readreg_25(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[25]~q ),
	.break_readreg_5(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[5]~q ),
	.jdo_7(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[7]~q ),
	.jdo_24(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[24]~q ),
	.break_readreg_18(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[18]~q ),
	.break_readreg_21(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[21]~q ),
	.jdo_22(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[22]~q ),
	.jdo_14(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[14]~q ),
	.jdo_15(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[15]~q ),
	.jdo_8(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[8]~q ),
	.jdo_13(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[13]~q ),
	.jdo_12(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[12]~q ),
	.jdo_11(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[11]~q ),
	.jdo_10(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[10]~q ),
	.jdo_9(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[9]~q ),
	.break_readreg_6(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[6]~q ),
	.break_readreg_22(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[22]~q ),
	.break_readreg_15(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[15]~q ),
	.break_readreg_7(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[7]~q ),
	.break_readreg_23(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[23]~q ),
	.break_readreg_13(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[13]~q ),
	.break_readreg_14(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[14]~q ),
	.break_readreg_12(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[12]~q ),
	.break_readreg_11(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[11]~q ),
	.break_readreg_10(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[10]~q ),
	.break_readreg_9(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[9]~q ),
	.break_readreg_8(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[8]~q ),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3),
	.irf_reg_0_2(irf_reg_0_2),
	.irf_reg_1_2(irf_reg_1_2),
	.clk_clk(clk_clk));

nios_mcu_nios_mcu_nios_cpu_cpu_nios2_ocimem the_nios_mcu_nios_cpu_cpu_nios2_ocimem(
	.q_a_0(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[0] ),
	.q_a_1(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[1] ),
	.q_a_2(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[2] ),
	.q_a_22(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[22] ),
	.q_a_23(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[23] ),
	.q_a_24(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[24] ),
	.q_a_25(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[25] ),
	.q_a_26(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[26] ),
	.q_a_11(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[11] ),
	.q_a_13(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[13] ),
	.q_a_16(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[16] ),
	.q_a_12(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[12] ),
	.q_a_3(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[3] ),
	.q_a_5(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[5] ),
	.q_a_4(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[4] ),
	.q_a_14(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[14] ),
	.q_a_15(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[15] ),
	.q_a_18(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[18] ),
	.q_a_17(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[17] ),
	.q_a_10(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[10] ),
	.q_a_9(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[9] ),
	.q_a_8(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[8] ),
	.q_a_7(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[7] ),
	.q_a_6(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[6] ),
	.q_a_21(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[21] ),
	.q_a_19(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[19] ),
	.q_a_20(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[20] ),
	.MonDReg_4(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[4]~q ),
	.MonDReg_12(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[12]~q ),
	.MonDReg_5(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[5]~q ),
	.MonDReg_18(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[18]~q ),
	.q_a_27(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[27] ),
	.q_a_28(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[28] ),
	.q_a_29(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[29] ),
	.q_a_30(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[30] ),
	.q_a_31(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[31] ),
	.MonDReg_8(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[8]~q ),
	.MonDReg_29(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[29]~q ),
	.waitrequest1(waitrequest),
	.MonDReg_0(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[0]~q ),
	.write(\write~q ),
	.address_8(\address[8]~q ),
	.read(\read~q ),
	.MonDReg_1(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[1]~q ),
	.jdo_3(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[3]~q ),
	.jdo_35(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[35]~q ),
	.take_action_ocimem_b(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|take_action_ocimem_b~combout ),
	.take_action_ocimem_a(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~0_combout ),
	.jdo_17(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[17]~q ),
	.take_action_ocimem_a1(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~1_combout ),
	.jdo_34(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[34]~q ),
	.MonDReg_2(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[2]~q ),
	.jdo_4(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[4]~q ),
	.debugaccess(\debugaccess~q ),
	.r_early_rst(r_early_rst),
	.writedata_0(\writedata[0]~q ),
	.address_0(\address[0]~q ),
	.address_1(\address[1]~q ),
	.address_2(\address[2]~q ),
	.address_3(\address[3]~q ),
	.address_4(\address[4]~q ),
	.address_5(\address[5]~q ),
	.address_6(\address[6]~q ),
	.address_7(\address[7]~q ),
	.byteenable_0(\byteenable[0]~q ),
	.jdo_25(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[25]~q ),
	.jdo_21(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[21]~q ),
	.jdo_20(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[20]~q ),
	.jdo_33(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[33]~q ),
	.jdo_32(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[32]~q ),
	.jdo_31(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[31]~q ),
	.jdo_30(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[30]~q ),
	.jdo_29(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[29]~q ),
	.jdo_28(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[28]~q ),
	.jdo_27(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[27]~q ),
	.jdo_26(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[26]~q ),
	.MonDReg_3(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[3]~q ),
	.jdo_5(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[5]~q ),
	.writedata_1(\writedata[1]~q ),
	.jdo_19(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[19]~q ),
	.jdo_18(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[18]~q ),
	.writedata_3(\writedata[3]~q ),
	.MonDReg_16(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[16]~q ),
	.jdo_6(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[6]~q ),
	.writedata_2(\writedata[2]~q ),
	.MonDReg_24(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[24]~q ),
	.MonDReg_20(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[20]~q ),
	.MonDReg_19(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[19]~q ),
	.MonDReg_22(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[22]~q ),
	.writedata_22(\writedata[22]~q ),
	.byteenable_2(\byteenable[2]~q ),
	.MonDReg_23(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[23]~q ),
	.writedata_23(\writedata[23]~q ),
	.writedata_24(\writedata[24]~q ),
	.byteenable_3(\byteenable[3]~q ),
	.MonDReg_25(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[25]~q ),
	.writedata_25(\writedata[25]~q ),
	.MonDReg_26(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[26]~q ),
	.writedata_26(\writedata[26]~q ),
	.MonDReg_11(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[11]~q ),
	.writedata_11(\writedata[11]~q ),
	.byteenable_1(\byteenable[1]~q ),
	.MonDReg_13(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[13]~q ),
	.writedata_13(\writedata[13]~q ),
	.writedata_16(\writedata[16]~q ),
	.writedata_12(\writedata[12]~q ),
	.jdo_23(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[23]~q ),
	.writedata_5(\writedata[5]~q ),
	.writedata_4(\writedata[4]~q ),
	.MonDReg_14(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[14]~q ),
	.writedata_14(\writedata[14]~q ),
	.MonDReg_15(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[15]~q ),
	.writedata_15(\writedata[15]~q ),
	.writedata_18(\writedata[18]~q ),
	.MonDReg_17(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[17]~q ),
	.writedata_17(\writedata[17]~q ),
	.MonDReg_10(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[10]~q ),
	.writedata_10(\writedata[10]~q ),
	.MonDReg_9(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[9]~q ),
	.writedata_9(\writedata[9]~q ),
	.writedata_8(\writedata[8]~q ),
	.MonDReg_7(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[7]~q ),
	.writedata_7(\writedata[7]~q ),
	.MonDReg_6(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[6]~q ),
	.writedata_6(\writedata[6]~q ),
	.MonDReg_21(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[21]~q ),
	.writedata_21(\writedata[21]~q ),
	.writedata_19(\writedata[19]~q ),
	.writedata_20(\writedata[20]~q ),
	.jdo_16(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[16]~q ),
	.MonDReg_31(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[31]~q ),
	.MonDReg_30(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[30]~q ),
	.MonDReg_28(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[28]~q ),
	.MonDReg_27(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|MonDReg[27]~q ),
	.jdo_7(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[7]~q ),
	.jdo_24(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[24]~q ),
	.jdo_22(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[22]~q ),
	.jdo_14(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[14]~q ),
	.jdo_15(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[15]~q ),
	.jdo_8(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[8]~q ),
	.writedata_27(\writedata[27]~q ),
	.writedata_28(\writedata[28]~q ),
	.writedata_29(\writedata[29]~q ),
	.writedata_30(\writedata[30]~q ),
	.writedata_31(\writedata[31]~q ),
	.jdo_13(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[13]~q ),
	.jdo_12(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[12]~q ),
	.jdo_11(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[11]~q ),
	.jdo_10(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[10]~q ),
	.jdo_9(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[9]~q ),
	.clk_clk(clk_clk));

nios_mcu_nios_mcu_nios_cpu_cpu_nios2_avalon_reg the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg(
	.r_sync_rst(r_sync_rst),
	.write(\write~q ),
	.address_8(\address[8]~q ),
	.debugaccess(\debugaccess~q ),
	.writedata_0(\writedata[0]~q ),
	.address_0(\address[0]~q ),
	.address_1(\address[1]~q ),
	.address_2(\address[2]~q ),
	.address_3(\address[3]~q ),
	.address_4(\address[4]~q ),
	.address_5(\address[5]~q ),
	.address_6(\address[6]~q ),
	.address_7(\address[7]~q ),
	.Equal0(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|Equal0~2_combout ),
	.take_action_ocireg(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|take_action_ocireg~0_combout ),
	.oci_ienable_0(oci_ienable_0),
	.oci_single_step_mode1(oci_single_step_mode),
	.monitor_error(\the_nios_mcu_nios_cpu_cpu_nios2_oci_debug|monitor_error~q ),
	.Equal1(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.oci_reg_readdata_0(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_reg_readdata[0]~0_combout ),
	.writedata_3(\writedata[3]~q ),
	.oci_ienable_16(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.clk_clk(clk_clk));

nios_mcu_nios_mcu_nios_cpu_cpu_nios2_oci_break the_nios_mcu_nios_cpu_cpu_nios2_oci_break(
	.break_readreg_0(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[0]~q ),
	.break_readreg_1(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[1]~q ),
	.jdo_0(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[0]~q ),
	.jdo_36(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[36]~q ),
	.jdo_37(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[37]~q ),
	.ir_0(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|ir[0]~q ),
	.ir_1(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|ir[1]~q ),
	.enable_action_strobe(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|enable_action_strobe~q ),
	.jdo_3(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[3]~q ),
	.jdo_17(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[17]~q ),
	.break_readreg_2(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[2]~q ),
	.jdo_1(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[1]~q ),
	.jdo_4(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[4]~q ),
	.jdo_25(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[25]~q ),
	.jdo_21(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[21]~q ),
	.jdo_20(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[20]~q ),
	.jdo_31(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[31]~q ),
	.jdo_30(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[30]~q ),
	.jdo_29(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[29]~q ),
	.jdo_28(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[28]~q ),
	.jdo_27(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[27]~q ),
	.jdo_26(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[26]~q ),
	.break_readreg_3(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[3]~q ),
	.jdo_2(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[2]~q ),
	.jdo_5(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[5]~q ),
	.jdo_19(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[19]~q ),
	.jdo_18(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[18]~q ),
	.break_readreg_16(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[16]~q ),
	.break_readreg_4(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[4]~q ),
	.jdo_6(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[6]~q ),
	.break_readreg_24(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[24]~q ),
	.break_readreg_20(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[20]~q ),
	.break_readreg_19(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[19]~q ),
	.jdo_23(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[23]~q ),
	.break_readreg_17(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[17]~q ),
	.jdo_16(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[16]~q ),
	.break_readreg_31(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[31]~q ),
	.break_readreg_30(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[30]~q ),
	.break_readreg_29(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[29]~q ),
	.break_readreg_28(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[28]~q ),
	.break_readreg_27(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[27]~q ),
	.break_readreg_26(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[26]~q ),
	.break_readreg_25(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[25]~q ),
	.break_readreg_5(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[5]~q ),
	.jdo_7(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[7]~q ),
	.jdo_24(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[24]~q ),
	.break_readreg_18(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[18]~q ),
	.break_readreg_21(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[21]~q ),
	.jdo_22(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[22]~q ),
	.jdo_14(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[14]~q ),
	.jdo_15(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[15]~q ),
	.jdo_8(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[8]~q ),
	.jdo_13(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[13]~q ),
	.jdo_12(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[12]~q ),
	.jdo_11(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[11]~q ),
	.jdo_10(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[10]~q ),
	.jdo_9(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[9]~q ),
	.break_readreg_6(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[6]~q ),
	.break_readreg_22(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[22]~q ),
	.break_readreg_15(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[15]~q ),
	.break_readreg_7(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[7]~q ),
	.break_readreg_23(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[23]~q ),
	.break_readreg_13(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[13]~q ),
	.break_readreg_14(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[14]~q ),
	.break_readreg_12(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[12]~q ),
	.break_readreg_11(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[11]~q ),
	.break_readreg_10(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[10]~q ),
	.break_readreg_9(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[9]~q ),
	.break_readreg_8(\the_nios_mcu_nios_cpu_cpu_nios2_oci_break|break_readreg[8]~q ),
	.clk_clk(clk_clk));

nios_mcu_nios_mcu_nios_cpu_cpu_nios2_oci_debug the_nios_mcu_nios_cpu_cpu_nios2_oci_debug(
	.jtag_break1(jtag_break),
	.r_sync_rst(r_sync_rst),
	.monitor_ready1(\the_nios_mcu_nios_cpu_cpu_nios2_oci_debug|monitor_ready~q ),
	.take_action_ocimem_a(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~1_combout ),
	.jdo_34(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[34]~q ),
	.writedata_0(\writedata[0]~q ),
	.take_action_ocireg(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|take_action_ocireg~0_combout ),
	.jdo_25(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[25]~q ),
	.jdo_21(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[21]~q ),
	.jdo_20(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[20]~q ),
	.take_action_ocimem_a1(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|take_action_ocimem_a~combout ),
	.writedata_1(\writedata[1]~q ),
	.monitor_error1(\the_nios_mcu_nios_cpu_cpu_nios2_oci_debug|monitor_error~q ),
	.jdo_19(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[19]~q ),
	.jdo_18(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[18]~q ),
	.monitor_go1(\the_nios_mcu_nios_cpu_cpu_nios2_oci_debug|monitor_go~q ),
	.jdo_23(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[23]~q ),
	.resetlatch1(\the_nios_mcu_nios_cpu_cpu_nios2_oci_debug|resetlatch~q ),
	.jdo_24(\the_nios_mcu_nios_cpu_cpu_debug_slave_wrapper|the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk|jdo[24]~q ),
	.state_1(state_1),
	.clk_clk(clk_clk));

dffeas write(
	.clk(clk_clk),
	.d(\write~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\write~q ),
	.prn(vcc));
defparam write.is_wysiwyg = "true";
defparam write.power_up = "low";

dffeas read(
	.clk(clk_clk),
	.d(\read~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read~q ),
	.prn(vcc));
defparam read.is_wysiwyg = "true";
defparam read.power_up = "low";

cycloneive_lcell_comb \write~0 (
	.dataa(m0_write),
	.datab(saved_grant_0),
	.datac(mem_used_1),
	.datad(\write~q ),
	.cin(gnd),
	.combout(\write~0_combout ),
	.cout());
defparam \write~0 .lut_mask = 16'hEFFF;
defparam \write~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \write~1 (
	.dataa(waitrequest),
	.datab(WideOr1),
	.datac(\write~0_combout ),
	.datad(\write~q ),
	.cin(gnd),
	.combout(\write~1_combout ),
	.cout());
defparam \write~1 .lut_mask = 16'hFFFE;
defparam \write~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read~0 (
	.dataa(waitrequest),
	.datab(\read~q ),
	.datac(rf_source_valid),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\read~0_combout ),
	.cout());
defparam \read~0 .lut_mask = 16'hB8FF;
defparam \read~0 .sum_lutc_input = "datac";

dffeas debugaccess(
	.clk(clk_clk),
	.d(debugaccess_nxt),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\debugaccess~q ),
	.prn(vcc));
defparam debugaccess.is_wysiwyg = "true";
defparam debugaccess.power_up = "low";

dffeas \writedata[0] (
	.clk(clk_clk),
	.d(writedata_nxt[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[0]~q ),
	.prn(vcc));
defparam \writedata[0] .is_wysiwyg = "true";
defparam \writedata[0] .power_up = "low";

dffeas \address[0] (
	.clk(clk_clk),
	.d(address_nxt[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[0]~q ),
	.prn(vcc));
defparam \address[0] .is_wysiwyg = "true";
defparam \address[0] .power_up = "low";

dffeas \address[1] (
	.clk(clk_clk),
	.d(address_nxt[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[1]~q ),
	.prn(vcc));
defparam \address[1] .is_wysiwyg = "true";
defparam \address[1] .power_up = "low";

dffeas \address[2] (
	.clk(clk_clk),
	.d(address_nxt[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[2]~q ),
	.prn(vcc));
defparam \address[2] .is_wysiwyg = "true";
defparam \address[2] .power_up = "low";

dffeas \address[3] (
	.clk(clk_clk),
	.d(address_nxt[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[3]~q ),
	.prn(vcc));
defparam \address[3] .is_wysiwyg = "true";
defparam \address[3] .power_up = "low";

dffeas \address[4] (
	.clk(clk_clk),
	.d(address_nxt[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[4]~q ),
	.prn(vcc));
defparam \address[4] .is_wysiwyg = "true";
defparam \address[4] .power_up = "low";

dffeas \address[5] (
	.clk(clk_clk),
	.d(address_nxt[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[5]~q ),
	.prn(vcc));
defparam \address[5] .is_wysiwyg = "true";
defparam \address[5] .power_up = "low";

dffeas \address[6] (
	.clk(clk_clk),
	.d(address_nxt[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[6]~q ),
	.prn(vcc));
defparam \address[6] .is_wysiwyg = "true";
defparam \address[6] .power_up = "low";

dffeas \address[7] (
	.clk(clk_clk),
	.d(address_nxt[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[7]~q ),
	.prn(vcc));
defparam \address[7] .is_wysiwyg = "true";
defparam \address[7] .power_up = "low";

dffeas \byteenable[0] (
	.clk(clk_clk),
	.d(byteenable_nxt[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[0]~q ),
	.prn(vcc));
defparam \byteenable[0] .is_wysiwyg = "true";
defparam \byteenable[0] .power_up = "low";

dffeas \writedata[1] (
	.clk(clk_clk),
	.d(writedata_nxt[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[1]~q ),
	.prn(vcc));
defparam \writedata[1] .is_wysiwyg = "true";
defparam \writedata[1] .power_up = "low";

dffeas \writedata[3] (
	.clk(clk_clk),
	.d(writedata_nxt[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[3]~q ),
	.prn(vcc));
defparam \writedata[3] .is_wysiwyg = "true";
defparam \writedata[3] .power_up = "low";

dffeas \writedata[2] (
	.clk(clk_clk),
	.d(writedata_nxt[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[2]~q ),
	.prn(vcc));
defparam \writedata[2] .is_wysiwyg = "true";
defparam \writedata[2] .power_up = "low";

dffeas \writedata[22] (
	.clk(clk_clk),
	.d(writedata_nxt[22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[22]~q ),
	.prn(vcc));
defparam \writedata[22] .is_wysiwyg = "true";
defparam \writedata[22] .power_up = "low";

dffeas \byteenable[2] (
	.clk(clk_clk),
	.d(byteenable_nxt[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[2]~q ),
	.prn(vcc));
defparam \byteenable[2] .is_wysiwyg = "true";
defparam \byteenable[2] .power_up = "low";

dffeas \writedata[23] (
	.clk(clk_clk),
	.d(writedata_nxt[23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[23]~q ),
	.prn(vcc));
defparam \writedata[23] .is_wysiwyg = "true";
defparam \writedata[23] .power_up = "low";

dffeas \writedata[24] (
	.clk(clk_clk),
	.d(writedata_nxt[24]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[24]~q ),
	.prn(vcc));
defparam \writedata[24] .is_wysiwyg = "true";
defparam \writedata[24] .power_up = "low";

dffeas \byteenable[3] (
	.clk(clk_clk),
	.d(byteenable_nxt[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[3]~q ),
	.prn(vcc));
defparam \byteenable[3] .is_wysiwyg = "true";
defparam \byteenable[3] .power_up = "low";

dffeas \writedata[25] (
	.clk(clk_clk),
	.d(writedata_nxt[25]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[25]~q ),
	.prn(vcc));
defparam \writedata[25] .is_wysiwyg = "true";
defparam \writedata[25] .power_up = "low";

dffeas \writedata[26] (
	.clk(clk_clk),
	.d(writedata_nxt[26]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[26]~q ),
	.prn(vcc));
defparam \writedata[26] .is_wysiwyg = "true";
defparam \writedata[26] .power_up = "low";

dffeas \writedata[11] (
	.clk(clk_clk),
	.d(writedata_nxt[11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[11]~q ),
	.prn(vcc));
defparam \writedata[11] .is_wysiwyg = "true";
defparam \writedata[11] .power_up = "low";

dffeas \byteenable[1] (
	.clk(clk_clk),
	.d(byteenable_nxt[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[1]~q ),
	.prn(vcc));
defparam \byteenable[1] .is_wysiwyg = "true";
defparam \byteenable[1] .power_up = "low";

dffeas \writedata[13] (
	.clk(clk_clk),
	.d(writedata_nxt[13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[13]~q ),
	.prn(vcc));
defparam \writedata[13] .is_wysiwyg = "true";
defparam \writedata[13] .power_up = "low";

dffeas \writedata[16] (
	.clk(clk_clk),
	.d(writedata_nxt[16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[16]~q ),
	.prn(vcc));
defparam \writedata[16] .is_wysiwyg = "true";
defparam \writedata[16] .power_up = "low";

dffeas \writedata[12] (
	.clk(clk_clk),
	.d(writedata_nxt[12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[12]~q ),
	.prn(vcc));
defparam \writedata[12] .is_wysiwyg = "true";
defparam \writedata[12] .power_up = "low";

dffeas \writedata[5] (
	.clk(clk_clk),
	.d(writedata_nxt[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[5]~q ),
	.prn(vcc));
defparam \writedata[5] .is_wysiwyg = "true";
defparam \writedata[5] .power_up = "low";

dffeas \writedata[4] (
	.clk(clk_clk),
	.d(writedata_nxt[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[4]~q ),
	.prn(vcc));
defparam \writedata[4] .is_wysiwyg = "true";
defparam \writedata[4] .power_up = "low";

dffeas \writedata[14] (
	.clk(clk_clk),
	.d(writedata_nxt[14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[14]~q ),
	.prn(vcc));
defparam \writedata[14] .is_wysiwyg = "true";
defparam \writedata[14] .power_up = "low";

dffeas \writedata[15] (
	.clk(clk_clk),
	.d(writedata_nxt[15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[15]~q ),
	.prn(vcc));
defparam \writedata[15] .is_wysiwyg = "true";
defparam \writedata[15] .power_up = "low";

dffeas \writedata[18] (
	.clk(clk_clk),
	.d(writedata_nxt[18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[18]~q ),
	.prn(vcc));
defparam \writedata[18] .is_wysiwyg = "true";
defparam \writedata[18] .power_up = "low";

dffeas \writedata[17] (
	.clk(clk_clk),
	.d(writedata_nxt[17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[17]~q ),
	.prn(vcc));
defparam \writedata[17] .is_wysiwyg = "true";
defparam \writedata[17] .power_up = "low";

dffeas \writedata[10] (
	.clk(clk_clk),
	.d(writedata_nxt[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[10]~q ),
	.prn(vcc));
defparam \writedata[10] .is_wysiwyg = "true";
defparam \writedata[10] .power_up = "low";

dffeas \writedata[9] (
	.clk(clk_clk),
	.d(writedata_nxt[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[9]~q ),
	.prn(vcc));
defparam \writedata[9] .is_wysiwyg = "true";
defparam \writedata[9] .power_up = "low";

dffeas \writedata[8] (
	.clk(clk_clk),
	.d(writedata_nxt[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[8]~q ),
	.prn(vcc));
defparam \writedata[8] .is_wysiwyg = "true";
defparam \writedata[8] .power_up = "low";

dffeas \writedata[7] (
	.clk(clk_clk),
	.d(writedata_nxt[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[7]~q ),
	.prn(vcc));
defparam \writedata[7] .is_wysiwyg = "true";
defparam \writedata[7] .power_up = "low";

dffeas \writedata[6] (
	.clk(clk_clk),
	.d(writedata_nxt[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[6]~q ),
	.prn(vcc));
defparam \writedata[6] .is_wysiwyg = "true";
defparam \writedata[6] .power_up = "low";

dffeas \writedata[21] (
	.clk(clk_clk),
	.d(writedata_nxt[21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[21]~q ),
	.prn(vcc));
defparam \writedata[21] .is_wysiwyg = "true";
defparam \writedata[21] .power_up = "low";

dffeas \writedata[19] (
	.clk(clk_clk),
	.d(writedata_nxt[19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[19]~q ),
	.prn(vcc));
defparam \writedata[19] .is_wysiwyg = "true";
defparam \writedata[19] .power_up = "low";

dffeas \writedata[20] (
	.clk(clk_clk),
	.d(writedata_nxt[20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[20]~q ),
	.prn(vcc));
defparam \writedata[20] .is_wysiwyg = "true";
defparam \writedata[20] .power_up = "low";

dffeas \writedata[27] (
	.clk(clk_clk),
	.d(writedata_nxt[27]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[27]~q ),
	.prn(vcc));
defparam \writedata[27] .is_wysiwyg = "true";
defparam \writedata[27] .power_up = "low";

dffeas \writedata[28] (
	.clk(clk_clk),
	.d(writedata_nxt[28]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[28]~q ),
	.prn(vcc));
defparam \writedata[28] .is_wysiwyg = "true";
defparam \writedata[28] .power_up = "low";

dffeas \writedata[29] (
	.clk(clk_clk),
	.d(writedata_nxt[29]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[29]~q ),
	.prn(vcc));
defparam \writedata[29] .is_wysiwyg = "true";
defparam \writedata[29] .power_up = "low";

dffeas \writedata[30] (
	.clk(clk_clk),
	.d(writedata_nxt[30]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[30]~q ),
	.prn(vcc));
defparam \writedata[30] .is_wysiwyg = "true";
defparam \writedata[30] .power_up = "low";

dffeas \writedata[31] (
	.clk(clk_clk),
	.d(writedata_nxt[31]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[31]~q ),
	.prn(vcc));
defparam \writedata[31] .is_wysiwyg = "true";
defparam \writedata[31] .power_up = "low";

dffeas \readdata[0] (
	.clk(clk_clk),
	.d(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_reg_readdata[0]~0_combout ),
	.asdata(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[0] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas \readdata[1] (
	.clk(clk_clk),
	.d(\readdata~9_combout ),
	.asdata(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[1] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

dffeas \readdata[3] (
	.clk(clk_clk),
	.d(\readdata~10_combout ),
	.asdata(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[3] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_3),
	.prn(vcc));
defparam \readdata[3] .is_wysiwyg = "true";
defparam \readdata[3] .power_up = "low";

dffeas \readdata[2] (
	.clk(clk_clk),
	.d(\readdata~11_combout ),
	.asdata(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[2] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

dffeas \readdata[22] (
	.clk(clk_clk),
	.d(\readdata~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_22),
	.prn(vcc));
defparam \readdata[22] .is_wysiwyg = "true";
defparam \readdata[22] .power_up = "low";

dffeas \readdata[23] (
	.clk(clk_clk),
	.d(\readdata~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_23),
	.prn(vcc));
defparam \readdata[23] .is_wysiwyg = "true";
defparam \readdata[23] .power_up = "low";

dffeas \readdata[24] (
	.clk(clk_clk),
	.d(\readdata~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_24),
	.prn(vcc));
defparam \readdata[24] .is_wysiwyg = "true";
defparam \readdata[24] .power_up = "low";

dffeas \readdata[25] (
	.clk(clk_clk),
	.d(\readdata~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_25),
	.prn(vcc));
defparam \readdata[25] .is_wysiwyg = "true";
defparam \readdata[25] .power_up = "low";

dffeas \readdata[26] (
	.clk(clk_clk),
	.d(\readdata~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_26),
	.prn(vcc));
defparam \readdata[26] .is_wysiwyg = "true";
defparam \readdata[26] .power_up = "low";

dffeas \readdata[11] (
	.clk(clk_clk),
	.d(\readdata~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_11),
	.prn(vcc));
defparam \readdata[11] .is_wysiwyg = "true";
defparam \readdata[11] .power_up = "low";

dffeas \readdata[13] (
	.clk(clk_clk),
	.d(\readdata~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_13),
	.prn(vcc));
defparam \readdata[13] .is_wysiwyg = "true";
defparam \readdata[13] .power_up = "low";

dffeas \readdata[16] (
	.clk(clk_clk),
	.d(\readdata~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_16),
	.prn(vcc));
defparam \readdata[16] .is_wysiwyg = "true";
defparam \readdata[16] .power_up = "low";

dffeas \readdata[12] (
	.clk(clk_clk),
	.d(\readdata~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_12),
	.prn(vcc));
defparam \readdata[12] .is_wysiwyg = "true";
defparam \readdata[12] .power_up = "low";

dffeas \readdata[5] (
	.clk(clk_clk),
	.d(\readdata~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_5),
	.prn(vcc));
defparam \readdata[5] .is_wysiwyg = "true";
defparam \readdata[5] .power_up = "low";

dffeas \readdata[4] (
	.clk(clk_clk),
	.d(\readdata~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_4),
	.prn(vcc));
defparam \readdata[4] .is_wysiwyg = "true";
defparam \readdata[4] .power_up = "low";

dffeas \readdata[14] (
	.clk(clk_clk),
	.d(\readdata~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_14),
	.prn(vcc));
defparam \readdata[14] .is_wysiwyg = "true";
defparam \readdata[14] .power_up = "low";

dffeas \readdata[15] (
	.clk(clk_clk),
	.d(\readdata~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_15),
	.prn(vcc));
defparam \readdata[15] .is_wysiwyg = "true";
defparam \readdata[15] .power_up = "low";

dffeas \readdata[18] (
	.clk(clk_clk),
	.d(\readdata~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_18),
	.prn(vcc));
defparam \readdata[18] .is_wysiwyg = "true";
defparam \readdata[18] .power_up = "low";

dffeas \readdata[17] (
	.clk(clk_clk),
	.d(\readdata~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_17),
	.prn(vcc));
defparam \readdata[17] .is_wysiwyg = "true";
defparam \readdata[17] .power_up = "low";

dffeas \readdata[10] (
	.clk(clk_clk),
	.d(\readdata~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_10),
	.prn(vcc));
defparam \readdata[10] .is_wysiwyg = "true";
defparam \readdata[10] .power_up = "low";

dffeas \readdata[9] (
	.clk(clk_clk),
	.d(\readdata~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_9),
	.prn(vcc));
defparam \readdata[9] .is_wysiwyg = "true";
defparam \readdata[9] .power_up = "low";

dffeas \readdata[8] (
	.clk(clk_clk),
	.d(\readdata~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_8),
	.prn(vcc));
defparam \readdata[8] .is_wysiwyg = "true";
defparam \readdata[8] .power_up = "low";

dffeas \readdata[7] (
	.clk(clk_clk),
	.d(\readdata~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_7),
	.prn(vcc));
defparam \readdata[7] .is_wysiwyg = "true";
defparam \readdata[7] .power_up = "low";

dffeas \readdata[6] (
	.clk(clk_clk),
	.d(\readdata~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_6),
	.prn(vcc));
defparam \readdata[6] .is_wysiwyg = "true";
defparam \readdata[6] .power_up = "low";

dffeas \readdata[21] (
	.clk(clk_clk),
	.d(\readdata~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_21),
	.prn(vcc));
defparam \readdata[21] .is_wysiwyg = "true";
defparam \readdata[21] .power_up = "low";

dffeas \readdata[19] (
	.clk(clk_clk),
	.d(\readdata~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_19),
	.prn(vcc));
defparam \readdata[19] .is_wysiwyg = "true";
defparam \readdata[19] .power_up = "low";

dffeas \readdata[20] (
	.clk(clk_clk),
	.d(\readdata~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_20),
	.prn(vcc));
defparam \readdata[20] .is_wysiwyg = "true";
defparam \readdata[20] .power_up = "low";

dffeas \readdata[27] (
	.clk(clk_clk),
	.d(\readdata~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_27),
	.prn(vcc));
defparam \readdata[27] .is_wysiwyg = "true";
defparam \readdata[27] .power_up = "low";

dffeas \readdata[28] (
	.clk(clk_clk),
	.d(\readdata~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_28),
	.prn(vcc));
defparam \readdata[28] .is_wysiwyg = "true";
defparam \readdata[28] .power_up = "low";

dffeas \readdata[29] (
	.clk(clk_clk),
	.d(\readdata~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_29),
	.prn(vcc));
defparam \readdata[29] .is_wysiwyg = "true";
defparam \readdata[29] .power_up = "low";

dffeas \readdata[30] (
	.clk(clk_clk),
	.d(\readdata~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_30),
	.prn(vcc));
defparam \readdata[30] .is_wysiwyg = "true";
defparam \readdata[30] .power_up = "low";

dffeas \readdata[31] (
	.clk(clk_clk),
	.d(\readdata~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_31),
	.prn(vcc));
defparam \readdata[31] .is_wysiwyg = "true";
defparam \readdata[31] .power_up = "low";

dffeas \address[8] (
	.clk(clk_clk),
	.d(address_nxt[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[8]~q ),
	.prn(vcc));
defparam \address[8] .is_wysiwyg = "true";
defparam \address[8] .power_up = "low";

cycloneive_lcell_comb \readdata~9 (
	.dataa(\the_nios_mcu_nios_cpu_cpu_nios2_oci_debug|monitor_ready~q ),
	.datab(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datac(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datad(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|Equal0~2_combout ),
	.cin(gnd),
	.combout(\readdata~9_combout ),
	.cout());
defparam \readdata~9 .lut_mask = 16'hFAFC;
defparam \readdata~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~10 (
	.dataa(oci_single_step_mode),
	.datab(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datac(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datad(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|Equal0~2_combout ),
	.cin(gnd),
	.combout(\readdata~10_combout ),
	.cout());
defparam \readdata~10 .lut_mask = 16'hFAFC;
defparam \readdata~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~11 (
	.dataa(\the_nios_mcu_nios_cpu_cpu_nios2_oci_debug|monitor_go~q ),
	.datab(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datac(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datad(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|Equal0~2_combout ),
	.cin(gnd),
	.combout(\readdata~11_combout ),
	.cout());
defparam \readdata~11 .lut_mask = 16'hFAFC;
defparam \readdata~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~0 (
	.dataa(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[22] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~0_combout ),
	.cout());
defparam \readdata~0 .lut_mask = 16'hFAFC;
defparam \readdata~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~1 (
	.dataa(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[23] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~1_combout ),
	.cout());
defparam \readdata~1 .lut_mask = 16'hFAFC;
defparam \readdata~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~2 (
	.dataa(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[24] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~2_combout ),
	.cout());
defparam \readdata~2 .lut_mask = 16'hFAFC;
defparam \readdata~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~3 (
	.dataa(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[25] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~3_combout ),
	.cout());
defparam \readdata~3 .lut_mask = 16'hFAFC;
defparam \readdata~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~4 (
	.dataa(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[26] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~4_combout ),
	.cout());
defparam \readdata~4 .lut_mask = 16'hFAFC;
defparam \readdata~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~5 (
	.dataa(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[11] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~5_combout ),
	.cout());
defparam \readdata~5 .lut_mask = 16'hFAFC;
defparam \readdata~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~6 (
	.dataa(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[13] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~6_combout ),
	.cout());
defparam \readdata~6 .lut_mask = 16'hFAFC;
defparam \readdata~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~7 (
	.dataa(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[16] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~7_combout ),
	.cout());
defparam \readdata~7 .lut_mask = 16'hFAFC;
defparam \readdata~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~8 (
	.dataa(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[12] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~8_combout ),
	.cout());
defparam \readdata~8 .lut_mask = 16'hFAFC;
defparam \readdata~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~12 (
	.dataa(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[5] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~12_combout ),
	.cout());
defparam \readdata~12 .lut_mask = 16'hFAFC;
defparam \readdata~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~13 (
	.dataa(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[4] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~13_combout ),
	.cout());
defparam \readdata~13 .lut_mask = 16'hFAFC;
defparam \readdata~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~14 (
	.dataa(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[14] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~14_combout ),
	.cout());
defparam \readdata~14 .lut_mask = 16'hFAFC;
defparam \readdata~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~15 (
	.dataa(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[15] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~15_combout ),
	.cout());
defparam \readdata~15 .lut_mask = 16'hFAFC;
defparam \readdata~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~16 (
	.dataa(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[18] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~16_combout ),
	.cout());
defparam \readdata~16 .lut_mask = 16'hFAFC;
defparam \readdata~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~17 (
	.dataa(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[17] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~17_combout ),
	.cout());
defparam \readdata~17 .lut_mask = 16'hFAFC;
defparam \readdata~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~18 (
	.dataa(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[10] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~18_combout ),
	.cout());
defparam \readdata~18 .lut_mask = 16'hFAFC;
defparam \readdata~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~19 (
	.dataa(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[9] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~19_combout ),
	.cout());
defparam \readdata~19 .lut_mask = 16'hFAFC;
defparam \readdata~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~20 (
	.dataa(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[8] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~20_combout ),
	.cout());
defparam \readdata~20 .lut_mask = 16'hFAFC;
defparam \readdata~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~21 (
	.dataa(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[7] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~21_combout ),
	.cout());
defparam \readdata~21 .lut_mask = 16'hFAFC;
defparam \readdata~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~22 (
	.dataa(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[6] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~22_combout ),
	.cout());
defparam \readdata~22 .lut_mask = 16'hFAFC;
defparam \readdata~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~23 (
	.dataa(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[21] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~23_combout ),
	.cout());
defparam \readdata~23 .lut_mask = 16'hFAFC;
defparam \readdata~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~24 (
	.dataa(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[19] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~24_combout ),
	.cout());
defparam \readdata~24 .lut_mask = 16'hFAFC;
defparam \readdata~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~25 (
	.dataa(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[20] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~25_combout ),
	.cout());
defparam \readdata~25 .lut_mask = 16'hFAFC;
defparam \readdata~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~26 (
	.dataa(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[27] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~26_combout ),
	.cout());
defparam \readdata~26 .lut_mask = 16'hFAFC;
defparam \readdata~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~27 (
	.dataa(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[28] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~27_combout ),
	.cout());
defparam \readdata~27 .lut_mask = 16'hFAFC;
defparam \readdata~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~28 (
	.dataa(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[29] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~28_combout ),
	.cout());
defparam \readdata~28 .lut_mask = 16'hFAFC;
defparam \readdata~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~29 (
	.dataa(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[30] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~29_combout ),
	.cout());
defparam \readdata~29 .lut_mask = 16'hFAFC;
defparam \readdata~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata~30 (
	.dataa(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datab(\the_nios_mcu_nios_cpu_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(\the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[31] ),
	.datad(\address[8]~q ),
	.cin(gnd),
	.combout(\readdata~30_combout ),
	.cout());
defparam \readdata~30 .lut_mask = 16'hFAFC;
defparam \readdata~30 .sum_lutc_input = "datac";

endmodule

module nios_mcu_nios_mcu_nios_cpu_cpu_debug_slave_wrapper (
	sr_0,
	MonDReg_4,
	MonDReg_12,
	MonDReg_5,
	MonDReg_18,
	MonDReg_8,
	MonDReg_29,
	ir_out_0,
	ir_out_1,
	break_readreg_0,
	MonDReg_0,
	break_readreg_1,
	MonDReg_1,
	jdo_0,
	jdo_36,
	jdo_37,
	ir_0,
	ir_1,
	enable_action_strobe,
	jdo_3,
	jdo_35,
	take_action_ocimem_b,
	take_action_ocimem_a,
	monitor_ready,
	hbreak_enabled,
	jdo_17,
	take_action_ocimem_a1,
	jdo_34,
	break_readreg_2,
	MonDReg_2,
	jdo_1,
	jdo_4,
	jdo_25,
	jdo_21,
	jdo_20,
	take_action_ocimem_a2,
	jdo_33,
	jdo_32,
	jdo_31,
	jdo_30,
	jdo_29,
	jdo_28,
	jdo_27,
	jdo_26,
	break_readreg_3,
	MonDReg_3,
	jdo_2,
	jdo_5,
	monitor_error,
	jdo_19,
	jdo_18,
	break_readreg_16,
	MonDReg_16,
	break_readreg_4,
	jdo_6,
	break_readreg_24,
	MonDReg_24,
	break_readreg_20,
	MonDReg_20,
	break_readreg_19,
	MonDReg_19,
	MonDReg_22,
	MonDReg_23,
	MonDReg_25,
	MonDReg_26,
	MonDReg_11,
	MonDReg_13,
	jdo_23,
	MonDReg_14,
	MonDReg_15,
	MonDReg_17,
	MonDReg_10,
	MonDReg_9,
	MonDReg_7,
	MonDReg_6,
	MonDReg_21,
	break_readreg_17,
	jdo_16,
	resetlatch,
	break_readreg_31,
	MonDReg_31,
	break_readreg_30,
	MonDReg_30,
	break_readreg_29,
	break_readreg_28,
	MonDReg_28,
	break_readreg_27,
	MonDReg_27,
	break_readreg_26,
	break_readreg_25,
	break_readreg_5,
	jdo_7,
	jdo_24,
	break_readreg_18,
	break_readreg_21,
	jdo_22,
	jdo_14,
	jdo_15,
	jdo_8,
	jdo_13,
	jdo_12,
	jdo_11,
	jdo_10,
	jdo_9,
	break_readreg_6,
	break_readreg_22,
	break_readreg_15,
	break_readreg_7,
	break_readreg_23,
	break_readreg_13,
	break_readreg_14,
	break_readreg_12,
	break_readreg_11,
	break_readreg_10,
	break_readreg_9,
	break_readreg_8,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	sr_0;
input 	MonDReg_4;
input 	MonDReg_12;
input 	MonDReg_5;
input 	MonDReg_18;
input 	MonDReg_8;
input 	MonDReg_29;
output 	ir_out_0;
output 	ir_out_1;
input 	break_readreg_0;
input 	MonDReg_0;
input 	break_readreg_1;
input 	MonDReg_1;
output 	jdo_0;
output 	jdo_36;
output 	jdo_37;
output 	ir_0;
output 	ir_1;
output 	enable_action_strobe;
output 	jdo_3;
output 	jdo_35;
output 	take_action_ocimem_b;
output 	take_action_ocimem_a;
input 	monitor_ready;
input 	hbreak_enabled;
output 	jdo_17;
output 	take_action_ocimem_a1;
output 	jdo_34;
input 	break_readreg_2;
input 	MonDReg_2;
output 	jdo_1;
output 	jdo_4;
output 	jdo_25;
output 	jdo_21;
output 	jdo_20;
output 	take_action_ocimem_a2;
output 	jdo_33;
output 	jdo_32;
output 	jdo_31;
output 	jdo_30;
output 	jdo_29;
output 	jdo_28;
output 	jdo_27;
output 	jdo_26;
input 	break_readreg_3;
input 	MonDReg_3;
output 	jdo_2;
output 	jdo_5;
input 	monitor_error;
output 	jdo_19;
output 	jdo_18;
input 	break_readreg_16;
input 	MonDReg_16;
input 	break_readreg_4;
output 	jdo_6;
input 	break_readreg_24;
input 	MonDReg_24;
input 	break_readreg_20;
input 	MonDReg_20;
input 	break_readreg_19;
input 	MonDReg_19;
input 	MonDReg_22;
input 	MonDReg_23;
input 	MonDReg_25;
input 	MonDReg_26;
input 	MonDReg_11;
input 	MonDReg_13;
output 	jdo_23;
input 	MonDReg_14;
input 	MonDReg_15;
input 	MonDReg_17;
input 	MonDReg_10;
input 	MonDReg_9;
input 	MonDReg_7;
input 	MonDReg_6;
input 	MonDReg_21;
input 	break_readreg_17;
output 	jdo_16;
input 	resetlatch;
input 	break_readreg_31;
input 	MonDReg_31;
input 	break_readreg_30;
input 	MonDReg_30;
input 	break_readreg_29;
input 	break_readreg_28;
input 	MonDReg_28;
input 	break_readreg_27;
input 	MonDReg_27;
input 	break_readreg_26;
input 	break_readreg_25;
input 	break_readreg_5;
output 	jdo_7;
output 	jdo_24;
input 	break_readreg_18;
input 	break_readreg_21;
output 	jdo_22;
output 	jdo_14;
output 	jdo_15;
output 	jdo_8;
output 	jdo_13;
output 	jdo_12;
output 	jdo_11;
output 	jdo_10;
output 	jdo_9;
input 	break_readreg_6;
input 	break_readreg_22;
input 	break_readreg_15;
input 	break_readreg_7;
input 	break_readreg_23;
input 	break_readreg_13;
input 	break_readreg_14;
input 	break_readreg_12;
input 	break_readreg_11;
input 	break_readreg_10;
input 	break_readreg_9;
input 	break_readreg_8;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[35]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[31]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[7]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[15]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[1]~q ;
wire \nios_mcu_nios_cpu_cpu_debug_slave_phy|virtual_state_cdr~combout ;
wire \nios_mcu_nios_cpu_cpu_debug_slave_phy|virtual_state_sdr~0_combout ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[2]~q ;
wire \nios_mcu_nios_cpu_cpu_debug_slave_phy|virtual_state_uir~0_combout ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[3]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[4]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[36]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[37]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[17]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[34]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[5]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[25]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[21]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[20]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[18]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[33]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[32]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[30]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[29]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[28]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[27]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[26]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[6]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[19]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[22]~q ;
wire \nios_mcu_nios_cpu_cpu_debug_slave_phy|virtual_state_udr~0_combout ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[23]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[16]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[8]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[24]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[14]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[13]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[12]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[11]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[10]~q ;
wire \the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[9]~q ;


nios_mcu_nios_mcu_nios_cpu_cpu_debug_slave_sysclk the_nios_mcu_nios_cpu_cpu_debug_slave_sysclk(
	.sr_0(sr_0),
	.sr_35(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[35]~q ),
	.sr_31(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[31]~q ),
	.sr_7(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[7]~q ),
	.sr_15(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[15]~q ),
	.sr_1(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[1]~q ),
	.sr_2(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[2]~q ),
	.virtual_state_uir(\nios_mcu_nios_cpu_cpu_debug_slave_phy|virtual_state_uir~0_combout ),
	.sr_3(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[3]~q ),
	.jdo_0(jdo_0),
	.jdo_36(jdo_36),
	.jdo_37(jdo_37),
	.ir_0(ir_0),
	.ir_1(ir_1),
	.enable_action_strobe1(enable_action_strobe),
	.jdo_3(jdo_3),
	.jdo_35(jdo_35),
	.take_action_ocimem_b1(take_action_ocimem_b),
	.take_action_ocimem_a1(take_action_ocimem_a),
	.jdo_17(jdo_17),
	.take_action_ocimem_a2(take_action_ocimem_a1),
	.jdo_34(jdo_34),
	.sr_4(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[4]~q ),
	.jdo_1(jdo_1),
	.jdo_4(jdo_4),
	.sr_36(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[36]~q ),
	.sr_37(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[37]~q ),
	.jdo_25(jdo_25),
	.jdo_21(jdo_21),
	.jdo_20(jdo_20),
	.take_action_ocimem_a3(take_action_ocimem_a2),
	.sr_17(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[17]~q ),
	.jdo_33(jdo_33),
	.jdo_32(jdo_32),
	.jdo_31(jdo_31),
	.jdo_30(jdo_30),
	.jdo_29(jdo_29),
	.jdo_28(jdo_28),
	.jdo_27(jdo_27),
	.jdo_26(jdo_26),
	.sr_34(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[34]~q ),
	.sr_5(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[5]~q ),
	.jdo_2(jdo_2),
	.jdo_5(jdo_5),
	.sr_25(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[25]~q ),
	.jdo_19(jdo_19),
	.jdo_18(jdo_18),
	.sr_21(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[21]~q ),
	.sr_20(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[20]~q ),
	.sr_18(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[18]~q ),
	.sr_33(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[33]~q ),
	.sr_32(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[32]~q ),
	.sr_30(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[30]~q ),
	.sr_29(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[29]~q ),
	.sr_28(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[28]~q ),
	.sr_27(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[27]~q ),
	.sr_26(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[26]~q ),
	.sr_6(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[6]~q ),
	.jdo_6(jdo_6),
	.sr_19(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[19]~q ),
	.sr_22(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[22]~q ),
	.jdo_23(jdo_23),
	.jdo_16(jdo_16),
	.jdo_7(jdo_7),
	.virtual_state_udr(\nios_mcu_nios_cpu_cpu_debug_slave_phy|virtual_state_udr~0_combout ),
	.jdo_24(jdo_24),
	.sr_23(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[23]~q ),
	.jdo_22(jdo_22),
	.jdo_14(jdo_14),
	.jdo_15(jdo_15),
	.jdo_8(jdo_8),
	.jdo_13(jdo_13),
	.jdo_12(jdo_12),
	.jdo_11(jdo_11),
	.jdo_10(jdo_10),
	.jdo_9(jdo_9),
	.sr_16(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[16]~q ),
	.sr_8(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[8]~q ),
	.sr_24(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[24]~q ),
	.sr_14(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[14]~q ),
	.sr_13(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[13]~q ),
	.sr_12(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[12]~q ),
	.sr_11(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[11]~q ),
	.sr_10(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[10]~q ),
	.sr_9(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[9]~q ),
	.ir_in({irf_reg_1_2,irf_reg_0_2}),
	.clk_clk(clk_clk));

nios_mcu_nios_mcu_nios_cpu_cpu_debug_slave_tck the_nios_mcu_nios_cpu_cpu_debug_slave_tck(
	.sr_0(sr_0),
	.sr_35(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[35]~q ),
	.sr_31(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[31]~q ),
	.MonDReg_4(MonDReg_4),
	.MonDReg_12(MonDReg_12),
	.MonDReg_5(MonDReg_5),
	.MonDReg_18(MonDReg_18),
	.MonDReg_8(MonDReg_8),
	.MonDReg_29(MonDReg_29),
	.sr_7(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[7]~q ),
	.sr_15(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[15]~q ),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.sr_1(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[1]~q ),
	.virtual_state_cdr(\nios_mcu_nios_cpu_cpu_debug_slave_phy|virtual_state_cdr~combout ),
	.virtual_state_sdr(\nios_mcu_nios_cpu_cpu_debug_slave_phy|virtual_state_sdr~0_combout ),
	.sr_2(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[2]~q ),
	.break_readreg_0(break_readreg_0),
	.MonDReg_0(MonDReg_0),
	.virtual_state_uir(\nios_mcu_nios_cpu_cpu_debug_slave_phy|virtual_state_uir~0_combout ),
	.sr_3(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[3]~q ),
	.break_readreg_1(break_readreg_1),
	.MonDReg_1(MonDReg_1),
	.monitor_ready(monitor_ready),
	.hbreak_enabled(hbreak_enabled),
	.sr_4(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[4]~q ),
	.break_readreg_2(break_readreg_2),
	.MonDReg_2(MonDReg_2),
	.sr_36(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[36]~q ),
	.sr_37(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[37]~q ),
	.sr_17(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[17]~q ),
	.sr_34(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[34]~q ),
	.sr_5(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[5]~q ),
	.break_readreg_3(break_readreg_3),
	.MonDReg_3(MonDReg_3),
	.sr_25(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[25]~q ),
	.monitor_error(monitor_error),
	.sr_21(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[21]~q ),
	.sr_20(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[20]~q ),
	.sr_18(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[18]~q ),
	.break_readreg_16(break_readreg_16),
	.MonDReg_16(MonDReg_16),
	.sr_33(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[33]~q ),
	.sr_32(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[32]~q ),
	.sr_30(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[30]~q ),
	.sr_29(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[29]~q ),
	.sr_28(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[28]~q ),
	.sr_27(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[27]~q ),
	.sr_26(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[26]~q ),
	.sr_6(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[6]~q ),
	.break_readreg_4(break_readreg_4),
	.break_readreg_24(break_readreg_24),
	.MonDReg_24(MonDReg_24),
	.sr_19(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[19]~q ),
	.sr_22(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[22]~q ),
	.break_readreg_20(break_readreg_20),
	.MonDReg_20(MonDReg_20),
	.break_readreg_19(break_readreg_19),
	.MonDReg_19(MonDReg_19),
	.MonDReg_22(MonDReg_22),
	.MonDReg_23(MonDReg_23),
	.MonDReg_25(MonDReg_25),
	.MonDReg_26(MonDReg_26),
	.MonDReg_11(MonDReg_11),
	.MonDReg_13(MonDReg_13),
	.MonDReg_14(MonDReg_14),
	.MonDReg_15(MonDReg_15),
	.MonDReg_17(MonDReg_17),
	.MonDReg_10(MonDReg_10),
	.MonDReg_9(MonDReg_9),
	.MonDReg_7(MonDReg_7),
	.MonDReg_6(MonDReg_6),
	.MonDReg_21(MonDReg_21),
	.break_readreg_17(break_readreg_17),
	.resetlatch(resetlatch),
	.break_readreg_31(break_readreg_31),
	.MonDReg_31(MonDReg_31),
	.break_readreg_30(break_readreg_30),
	.MonDReg_30(MonDReg_30),
	.break_readreg_29(break_readreg_29),
	.break_readreg_28(break_readreg_28),
	.MonDReg_28(MonDReg_28),
	.break_readreg_27(break_readreg_27),
	.MonDReg_27(MonDReg_27),
	.break_readreg_26(break_readreg_26),
	.break_readreg_25(break_readreg_25),
	.break_readreg_5(break_readreg_5),
	.break_readreg_18(break_readreg_18),
	.sr_23(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[23]~q ),
	.break_readreg_21(break_readreg_21),
	.sr_16(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[16]~q ),
	.break_readreg_6(break_readreg_6),
	.sr_8(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[8]~q ),
	.sr_24(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[24]~q ),
	.break_readreg_22(break_readreg_22),
	.sr_14(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[14]~q ),
	.sr_13(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[13]~q ),
	.sr_12(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[12]~q ),
	.sr_11(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[11]~q ),
	.sr_10(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[10]~q ),
	.sr_9(\the_nios_mcu_nios_cpu_cpu_debug_slave_tck|sr[9]~q ),
	.break_readreg_15(break_readreg_15),
	.break_readreg_7(break_readreg_7),
	.break_readreg_23(break_readreg_23),
	.break_readreg_13(break_readreg_13),
	.break_readreg_14(break_readreg_14),
	.break_readreg_12(break_readreg_12),
	.break_readreg_11(break_readreg_11),
	.break_readreg_10(break_readreg_10),
	.break_readreg_9(break_readreg_9),
	.break_readreg_8(break_readreg_8),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3),
	.irf_reg_0_2(irf_reg_0_2),
	.irf_reg_1_2(irf_reg_1_2));

nios_mcu_sld_virtual_jtag_basic_1 nios_mcu_nios_cpu_cpu_debug_slave_phy(
	.virtual_state_cdr1(\nios_mcu_nios_cpu_cpu_debug_slave_phy|virtual_state_cdr~combout ),
	.virtual_state_sdr(\nios_mcu_nios_cpu_cpu_debug_slave_phy|virtual_state_sdr~0_combout ),
	.virtual_state_uir(\nios_mcu_nios_cpu_cpu_debug_slave_phy|virtual_state_uir~0_combout ),
	.virtual_state_udr(\nios_mcu_nios_cpu_cpu_debug_slave_phy|virtual_state_udr~0_combout ),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3));

endmodule

module nios_mcu_nios_mcu_nios_cpu_cpu_debug_slave_sysclk (
	sr_0,
	sr_35,
	sr_31,
	sr_7,
	sr_15,
	sr_1,
	sr_2,
	virtual_state_uir,
	sr_3,
	jdo_0,
	jdo_36,
	jdo_37,
	ir_0,
	ir_1,
	enable_action_strobe1,
	jdo_3,
	jdo_35,
	take_action_ocimem_b1,
	take_action_ocimem_a1,
	jdo_17,
	take_action_ocimem_a2,
	jdo_34,
	sr_4,
	jdo_1,
	jdo_4,
	sr_36,
	sr_37,
	jdo_25,
	jdo_21,
	jdo_20,
	take_action_ocimem_a3,
	sr_17,
	jdo_33,
	jdo_32,
	jdo_31,
	jdo_30,
	jdo_29,
	jdo_28,
	jdo_27,
	jdo_26,
	sr_34,
	sr_5,
	jdo_2,
	jdo_5,
	sr_25,
	jdo_19,
	jdo_18,
	sr_21,
	sr_20,
	sr_18,
	sr_33,
	sr_32,
	sr_30,
	sr_29,
	sr_28,
	sr_27,
	sr_26,
	sr_6,
	jdo_6,
	sr_19,
	sr_22,
	jdo_23,
	jdo_16,
	jdo_7,
	virtual_state_udr,
	jdo_24,
	sr_23,
	jdo_22,
	jdo_14,
	jdo_15,
	jdo_8,
	jdo_13,
	jdo_12,
	jdo_11,
	jdo_10,
	jdo_9,
	sr_16,
	sr_8,
	sr_24,
	sr_14,
	sr_13,
	sr_12,
	sr_11,
	sr_10,
	sr_9,
	ir_in,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	sr_0;
input 	sr_35;
input 	sr_31;
input 	sr_7;
input 	sr_15;
input 	sr_1;
input 	sr_2;
input 	virtual_state_uir;
input 	sr_3;
output 	jdo_0;
output 	jdo_36;
output 	jdo_37;
output 	ir_0;
output 	ir_1;
output 	enable_action_strobe1;
output 	jdo_3;
output 	jdo_35;
output 	take_action_ocimem_b1;
output 	take_action_ocimem_a1;
output 	jdo_17;
output 	take_action_ocimem_a2;
output 	jdo_34;
input 	sr_4;
output 	jdo_1;
output 	jdo_4;
input 	sr_36;
input 	sr_37;
output 	jdo_25;
output 	jdo_21;
output 	jdo_20;
output 	take_action_ocimem_a3;
input 	sr_17;
output 	jdo_33;
output 	jdo_32;
output 	jdo_31;
output 	jdo_30;
output 	jdo_29;
output 	jdo_28;
output 	jdo_27;
output 	jdo_26;
input 	sr_34;
input 	sr_5;
output 	jdo_2;
output 	jdo_5;
input 	sr_25;
output 	jdo_19;
output 	jdo_18;
input 	sr_21;
input 	sr_20;
input 	sr_18;
input 	sr_33;
input 	sr_32;
input 	sr_30;
input 	sr_29;
input 	sr_28;
input 	sr_27;
input 	sr_26;
input 	sr_6;
output 	jdo_6;
input 	sr_19;
input 	sr_22;
output 	jdo_23;
output 	jdo_16;
output 	jdo_7;
input 	virtual_state_udr;
output 	jdo_24;
input 	sr_23;
output 	jdo_22;
output 	jdo_14;
output 	jdo_15;
output 	jdo_8;
output 	jdo_13;
output 	jdo_12;
output 	jdo_11;
output 	jdo_10;
output 	jdo_9;
input 	sr_16;
input 	sr_8;
input 	sr_24;
input 	sr_14;
input 	sr_13;
input 	sr_12;
input 	sr_11;
input 	sr_10;
input 	sr_9;
input 	[1:0] ir_in;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_altera_std_synchronizer3|dreg[0]~q ;
wire \the_altera_std_synchronizer4|dreg[0]~q ;
wire \sync2_udr~q ;
wire \update_jdo_strobe~0_combout ;
wire \update_jdo_strobe~q ;
wire \sync2_uir~q ;
wire \jxuir~0_combout ;
wire \jxuir~q ;


nios_mcu_altera_std_synchronizer_1 the_altera_std_synchronizer4(
	.din(virtual_state_uir),
	.dreg_0(\the_altera_std_synchronizer4|dreg[0]~q ),
	.clk(clk_clk));

nios_mcu_altera_std_synchronizer the_altera_std_synchronizer3(
	.dreg_0(\the_altera_std_synchronizer3|dreg[0]~q ),
	.din(virtual_state_udr),
	.clk(clk_clk));

dffeas \jdo[0] (
	.clk(clk_clk),
	.d(sr_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_0),
	.prn(vcc));
defparam \jdo[0] .is_wysiwyg = "true";
defparam \jdo[0] .power_up = "low";

dffeas \jdo[36] (
	.clk(clk_clk),
	.d(sr_36),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_36),
	.prn(vcc));
defparam \jdo[36] .is_wysiwyg = "true";
defparam \jdo[36] .power_up = "low";

dffeas \jdo[37] (
	.clk(clk_clk),
	.d(sr_37),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_37),
	.prn(vcc));
defparam \jdo[37] .is_wysiwyg = "true";
defparam \jdo[37] .power_up = "low";

dffeas \ir[0] (
	.clk(clk_clk),
	.d(ir_in[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\jxuir~q ),
	.q(ir_0),
	.prn(vcc));
defparam \ir[0] .is_wysiwyg = "true";
defparam \ir[0] .power_up = "low";

dffeas \ir[1] (
	.clk(clk_clk),
	.d(ir_in[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\jxuir~q ),
	.q(ir_1),
	.prn(vcc));
defparam \ir[1] .is_wysiwyg = "true";
defparam \ir[1] .power_up = "low";

dffeas enable_action_strobe(
	.clk(clk_clk),
	.d(\update_jdo_strobe~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(enable_action_strobe1),
	.prn(vcc));
defparam enable_action_strobe.is_wysiwyg = "true";
defparam enable_action_strobe.power_up = "low";

dffeas \jdo[3] (
	.clk(clk_clk),
	.d(sr_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_3),
	.prn(vcc));
defparam \jdo[3] .is_wysiwyg = "true";
defparam \jdo[3] .power_up = "low";

dffeas \jdo[35] (
	.clk(clk_clk),
	.d(sr_35),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_35),
	.prn(vcc));
defparam \jdo[35] .is_wysiwyg = "true";
defparam \jdo[35] .power_up = "low";

cycloneive_lcell_comb take_action_ocimem_b(
	.dataa(enable_action_strobe1),
	.datab(jdo_35),
	.datac(ir_1),
	.datad(ir_0),
	.cin(gnd),
	.combout(take_action_ocimem_b1),
	.cout());
defparam take_action_ocimem_b.lut_mask = 16'hEFFF;
defparam take_action_ocimem_b.sum_lutc_input = "datac";

cycloneive_lcell_comb \take_action_ocimem_a~0 (
	.dataa(enable_action_strobe1),
	.datab(gnd),
	.datac(ir_1),
	.datad(ir_0),
	.cin(gnd),
	.combout(take_action_ocimem_a1),
	.cout());
defparam \take_action_ocimem_a~0 .lut_mask = 16'hAFFF;
defparam \take_action_ocimem_a~0 .sum_lutc_input = "datac";

dffeas \jdo[17] (
	.clk(clk_clk),
	.d(sr_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_17),
	.prn(vcc));
defparam \jdo[17] .is_wysiwyg = "true";
defparam \jdo[17] .power_up = "low";

cycloneive_lcell_comb \take_action_ocimem_a~1 (
	.dataa(enable_action_strobe1),
	.datab(ir_1),
	.datac(ir_0),
	.datad(jdo_35),
	.cin(gnd),
	.combout(take_action_ocimem_a2),
	.cout());
defparam \take_action_ocimem_a~1 .lut_mask = 16'hBFFF;
defparam \take_action_ocimem_a~1 .sum_lutc_input = "datac";

dffeas \jdo[34] (
	.clk(clk_clk),
	.d(sr_34),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_34),
	.prn(vcc));
defparam \jdo[34] .is_wysiwyg = "true";
defparam \jdo[34] .power_up = "low";

dffeas \jdo[1] (
	.clk(clk_clk),
	.d(sr_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_1),
	.prn(vcc));
defparam \jdo[1] .is_wysiwyg = "true";
defparam \jdo[1] .power_up = "low";

dffeas \jdo[4] (
	.clk(clk_clk),
	.d(sr_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_4),
	.prn(vcc));
defparam \jdo[4] .is_wysiwyg = "true";
defparam \jdo[4] .power_up = "low";

dffeas \jdo[25] (
	.clk(clk_clk),
	.d(sr_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_25),
	.prn(vcc));
defparam \jdo[25] .is_wysiwyg = "true";
defparam \jdo[25] .power_up = "low";

dffeas \jdo[21] (
	.clk(clk_clk),
	.d(sr_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_21),
	.prn(vcc));
defparam \jdo[21] .is_wysiwyg = "true";
defparam \jdo[21] .power_up = "low";

dffeas \jdo[20] (
	.clk(clk_clk),
	.d(sr_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_20),
	.prn(vcc));
defparam \jdo[20] .is_wysiwyg = "true";
defparam \jdo[20] .power_up = "low";

cycloneive_lcell_comb take_action_ocimem_a(
	.dataa(take_action_ocimem_a1),
	.datab(jdo_34),
	.datac(gnd),
	.datad(jdo_35),
	.cin(gnd),
	.combout(take_action_ocimem_a3),
	.cout());
defparam take_action_ocimem_a.lut_mask = 16'hEEFF;
defparam take_action_ocimem_a.sum_lutc_input = "datac";

dffeas \jdo[33] (
	.clk(clk_clk),
	.d(sr_33),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_33),
	.prn(vcc));
defparam \jdo[33] .is_wysiwyg = "true";
defparam \jdo[33] .power_up = "low";

dffeas \jdo[32] (
	.clk(clk_clk),
	.d(sr_32),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_32),
	.prn(vcc));
defparam \jdo[32] .is_wysiwyg = "true";
defparam \jdo[32] .power_up = "low";

dffeas \jdo[31] (
	.clk(clk_clk),
	.d(sr_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_31),
	.prn(vcc));
defparam \jdo[31] .is_wysiwyg = "true";
defparam \jdo[31] .power_up = "low";

dffeas \jdo[30] (
	.clk(clk_clk),
	.d(sr_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_30),
	.prn(vcc));
defparam \jdo[30] .is_wysiwyg = "true";
defparam \jdo[30] .power_up = "low";

dffeas \jdo[29] (
	.clk(clk_clk),
	.d(sr_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_29),
	.prn(vcc));
defparam \jdo[29] .is_wysiwyg = "true";
defparam \jdo[29] .power_up = "low";

dffeas \jdo[28] (
	.clk(clk_clk),
	.d(sr_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_28),
	.prn(vcc));
defparam \jdo[28] .is_wysiwyg = "true";
defparam \jdo[28] .power_up = "low";

dffeas \jdo[27] (
	.clk(clk_clk),
	.d(sr_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_27),
	.prn(vcc));
defparam \jdo[27] .is_wysiwyg = "true";
defparam \jdo[27] .power_up = "low";

dffeas \jdo[26] (
	.clk(clk_clk),
	.d(sr_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_26),
	.prn(vcc));
defparam \jdo[26] .is_wysiwyg = "true";
defparam \jdo[26] .power_up = "low";

dffeas \jdo[2] (
	.clk(clk_clk),
	.d(sr_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_2),
	.prn(vcc));
defparam \jdo[2] .is_wysiwyg = "true";
defparam \jdo[2] .power_up = "low";

dffeas \jdo[5] (
	.clk(clk_clk),
	.d(sr_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_5),
	.prn(vcc));
defparam \jdo[5] .is_wysiwyg = "true";
defparam \jdo[5] .power_up = "low";

dffeas \jdo[19] (
	.clk(clk_clk),
	.d(sr_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_19),
	.prn(vcc));
defparam \jdo[19] .is_wysiwyg = "true";
defparam \jdo[19] .power_up = "low";

dffeas \jdo[18] (
	.clk(clk_clk),
	.d(sr_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_18),
	.prn(vcc));
defparam \jdo[18] .is_wysiwyg = "true";
defparam \jdo[18] .power_up = "low";

dffeas \jdo[6] (
	.clk(clk_clk),
	.d(sr_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_6),
	.prn(vcc));
defparam \jdo[6] .is_wysiwyg = "true";
defparam \jdo[6] .power_up = "low";

dffeas \jdo[23] (
	.clk(clk_clk),
	.d(sr_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_23),
	.prn(vcc));
defparam \jdo[23] .is_wysiwyg = "true";
defparam \jdo[23] .power_up = "low";

dffeas \jdo[16] (
	.clk(clk_clk),
	.d(sr_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_16),
	.prn(vcc));
defparam \jdo[16] .is_wysiwyg = "true";
defparam \jdo[16] .power_up = "low";

dffeas \jdo[7] (
	.clk(clk_clk),
	.d(sr_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_7),
	.prn(vcc));
defparam \jdo[7] .is_wysiwyg = "true";
defparam \jdo[7] .power_up = "low";

dffeas \jdo[24] (
	.clk(clk_clk),
	.d(sr_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_24),
	.prn(vcc));
defparam \jdo[24] .is_wysiwyg = "true";
defparam \jdo[24] .power_up = "low";

dffeas \jdo[22] (
	.clk(clk_clk),
	.d(sr_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_22),
	.prn(vcc));
defparam \jdo[22] .is_wysiwyg = "true";
defparam \jdo[22] .power_up = "low";

dffeas \jdo[14] (
	.clk(clk_clk),
	.d(sr_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_14),
	.prn(vcc));
defparam \jdo[14] .is_wysiwyg = "true";
defparam \jdo[14] .power_up = "low";

dffeas \jdo[15] (
	.clk(clk_clk),
	.d(sr_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_15),
	.prn(vcc));
defparam \jdo[15] .is_wysiwyg = "true";
defparam \jdo[15] .power_up = "low";

dffeas \jdo[8] (
	.clk(clk_clk),
	.d(sr_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_8),
	.prn(vcc));
defparam \jdo[8] .is_wysiwyg = "true";
defparam \jdo[8] .power_up = "low";

dffeas \jdo[13] (
	.clk(clk_clk),
	.d(sr_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_13),
	.prn(vcc));
defparam \jdo[13] .is_wysiwyg = "true";
defparam \jdo[13] .power_up = "low";

dffeas \jdo[12] (
	.clk(clk_clk),
	.d(sr_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_12),
	.prn(vcc));
defparam \jdo[12] .is_wysiwyg = "true";
defparam \jdo[12] .power_up = "low";

dffeas \jdo[11] (
	.clk(clk_clk),
	.d(sr_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_11),
	.prn(vcc));
defparam \jdo[11] .is_wysiwyg = "true";
defparam \jdo[11] .power_up = "low";

dffeas \jdo[10] (
	.clk(clk_clk),
	.d(sr_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_10),
	.prn(vcc));
defparam \jdo[10] .is_wysiwyg = "true";
defparam \jdo[10] .power_up = "low";

dffeas \jdo[9] (
	.clk(clk_clk),
	.d(sr_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_9),
	.prn(vcc));
defparam \jdo[9] .is_wysiwyg = "true";
defparam \jdo[9] .power_up = "low";

dffeas sync2_udr(
	.clk(clk_clk),
	.d(\the_altera_std_synchronizer3|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sync2_udr~q ),
	.prn(vcc));
defparam sync2_udr.is_wysiwyg = "true";
defparam sync2_udr.power_up = "low";

cycloneive_lcell_comb \update_jdo_strobe~0 (
	.dataa(\the_altera_std_synchronizer3|dreg[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\sync2_udr~q ),
	.cin(gnd),
	.combout(\update_jdo_strobe~0_combout ),
	.cout());
defparam \update_jdo_strobe~0 .lut_mask = 16'hAAFF;
defparam \update_jdo_strobe~0 .sum_lutc_input = "datac";

dffeas update_jdo_strobe(
	.clk(clk_clk),
	.d(\update_jdo_strobe~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\update_jdo_strobe~q ),
	.prn(vcc));
defparam update_jdo_strobe.is_wysiwyg = "true";
defparam update_jdo_strobe.power_up = "low";

dffeas sync2_uir(
	.clk(clk_clk),
	.d(\the_altera_std_synchronizer4|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sync2_uir~q ),
	.prn(vcc));
defparam sync2_uir.is_wysiwyg = "true";
defparam sync2_uir.power_up = "low";

cycloneive_lcell_comb \jxuir~0 (
	.dataa(\the_altera_std_synchronizer4|dreg[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\sync2_uir~q ),
	.cin(gnd),
	.combout(\jxuir~0_combout ),
	.cout());
defparam \jxuir~0 .lut_mask = 16'hAAFF;
defparam \jxuir~0 .sum_lutc_input = "datac";

dffeas jxuir(
	.clk(clk_clk),
	.d(\jxuir~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jxuir~q ),
	.prn(vcc));
defparam jxuir.is_wysiwyg = "true";
defparam jxuir.power_up = "low";

endmodule

module nios_mcu_altera_std_synchronizer (
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module nios_mcu_altera_std_synchronizer_1 (
	din,
	dreg_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	din;
output 	dreg_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module nios_mcu_nios_mcu_nios_cpu_cpu_debug_slave_tck (
	sr_0,
	sr_35,
	sr_31,
	MonDReg_4,
	MonDReg_12,
	MonDReg_5,
	MonDReg_18,
	MonDReg_8,
	MonDReg_29,
	sr_7,
	sr_15,
	ir_out_0,
	ir_out_1,
	sr_1,
	virtual_state_cdr,
	virtual_state_sdr,
	sr_2,
	break_readreg_0,
	MonDReg_0,
	virtual_state_uir,
	sr_3,
	break_readreg_1,
	MonDReg_1,
	monitor_ready,
	hbreak_enabled,
	sr_4,
	break_readreg_2,
	MonDReg_2,
	sr_36,
	sr_37,
	sr_17,
	sr_34,
	sr_5,
	break_readreg_3,
	MonDReg_3,
	sr_25,
	monitor_error,
	sr_21,
	sr_20,
	sr_18,
	break_readreg_16,
	MonDReg_16,
	sr_33,
	sr_32,
	sr_30,
	sr_29,
	sr_28,
	sr_27,
	sr_26,
	sr_6,
	break_readreg_4,
	break_readreg_24,
	MonDReg_24,
	sr_19,
	sr_22,
	break_readreg_20,
	MonDReg_20,
	break_readreg_19,
	MonDReg_19,
	MonDReg_22,
	MonDReg_23,
	MonDReg_25,
	MonDReg_26,
	MonDReg_11,
	MonDReg_13,
	MonDReg_14,
	MonDReg_15,
	MonDReg_17,
	MonDReg_10,
	MonDReg_9,
	MonDReg_7,
	MonDReg_6,
	MonDReg_21,
	break_readreg_17,
	resetlatch,
	break_readreg_31,
	MonDReg_31,
	break_readreg_30,
	MonDReg_30,
	break_readreg_29,
	break_readreg_28,
	MonDReg_28,
	break_readreg_27,
	MonDReg_27,
	break_readreg_26,
	break_readreg_25,
	break_readreg_5,
	break_readreg_18,
	sr_23,
	break_readreg_21,
	sr_16,
	break_readreg_6,
	sr_8,
	sr_24,
	break_readreg_22,
	sr_14,
	sr_13,
	sr_12,
	sr_11,
	sr_10,
	sr_9,
	break_readreg_15,
	break_readreg_7,
	break_readreg_23,
	break_readreg_13,
	break_readreg_14,
	break_readreg_12,
	break_readreg_11,
	break_readreg_10,
	break_readreg_9,
	break_readreg_8,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2)/* synthesis synthesis_greybox=1 */;
output 	sr_0;
output 	sr_35;
output 	sr_31;
input 	MonDReg_4;
input 	MonDReg_12;
input 	MonDReg_5;
input 	MonDReg_18;
input 	MonDReg_8;
input 	MonDReg_29;
output 	sr_7;
output 	sr_15;
output 	ir_out_0;
output 	ir_out_1;
output 	sr_1;
input 	virtual_state_cdr;
input 	virtual_state_sdr;
output 	sr_2;
input 	break_readreg_0;
input 	MonDReg_0;
input 	virtual_state_uir;
output 	sr_3;
input 	break_readreg_1;
input 	MonDReg_1;
input 	monitor_ready;
input 	hbreak_enabled;
output 	sr_4;
input 	break_readreg_2;
input 	MonDReg_2;
output 	sr_36;
output 	sr_37;
output 	sr_17;
output 	sr_34;
output 	sr_5;
input 	break_readreg_3;
input 	MonDReg_3;
output 	sr_25;
input 	monitor_error;
output 	sr_21;
output 	sr_20;
output 	sr_18;
input 	break_readreg_16;
input 	MonDReg_16;
output 	sr_33;
output 	sr_32;
output 	sr_30;
output 	sr_29;
output 	sr_28;
output 	sr_27;
output 	sr_26;
output 	sr_6;
input 	break_readreg_4;
input 	break_readreg_24;
input 	MonDReg_24;
output 	sr_19;
output 	sr_22;
input 	break_readreg_20;
input 	MonDReg_20;
input 	break_readreg_19;
input 	MonDReg_19;
input 	MonDReg_22;
input 	MonDReg_23;
input 	MonDReg_25;
input 	MonDReg_26;
input 	MonDReg_11;
input 	MonDReg_13;
input 	MonDReg_14;
input 	MonDReg_15;
input 	MonDReg_17;
input 	MonDReg_10;
input 	MonDReg_9;
input 	MonDReg_7;
input 	MonDReg_6;
input 	MonDReg_21;
input 	break_readreg_17;
input 	resetlatch;
input 	break_readreg_31;
input 	MonDReg_31;
input 	break_readreg_30;
input 	MonDReg_30;
input 	break_readreg_29;
input 	break_readreg_28;
input 	MonDReg_28;
input 	break_readreg_27;
input 	MonDReg_27;
input 	break_readreg_26;
input 	break_readreg_25;
input 	break_readreg_5;
input 	break_readreg_18;
output 	sr_23;
input 	break_readreg_21;
output 	sr_16;
input 	break_readreg_6;
output 	sr_8;
output 	sr_24;
input 	break_readreg_22;
output 	sr_14;
output 	sr_13;
output 	sr_12;
output 	sr_11;
output 	sr_10;
output 	sr_9;
input 	break_readreg_15;
input 	break_readreg_7;
input 	break_readreg_23;
input 	break_readreg_13;
input 	break_readreg_14;
input 	break_readreg_12;
input 	break_readreg_11;
input 	break_readreg_10;
input 	break_readreg_9;
input 	break_readreg_8;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_altera_std_synchronizer2|dreg[0]~q ;
wire \the_altera_std_synchronizer1|dreg[0]~q ;
wire \DRsize.000~q ;
wire \sr[0]~5_combout ;
wire \Mux37~0_combout ;
wire \sr~10_combout ;
wire \DRsize.100~q ;
wire \sr[35]~6_combout ;
wire \sr~23_combout ;
wire \sr~24_combout ;
wire \sr~25_combout ;
wire \sr[31]~44_combout ;
wire \sr[31]~7_combout ;
wire \Mux30~0_combout ;
wire \sr[7]~8_combout ;
wire \sr[33]~83_combout ;
wire \DRsize.010~q ;
wire \sr[15]~9_combout ;
wire \sr~71_combout ;
wire \sr~72_combout ;
wire \sr~11_combout ;
wire \sr~12_combout ;
wire \sr[14]~13_combout ;
wire \sr~14_combout ;
wire \sr~15_combout ;
wire \sr~16_combout ;
wire \sr~17_combout ;
wire \sr~18_combout ;
wire \sr~19_combout ;
wire \sr~20_combout ;
wire \sr[37]~21_combout ;
wire \sr~22_combout ;
wire \sr~26_combout ;
wire \sr~27_combout ;
wire \sr~28_combout ;
wire \sr[33]~29_combout ;
wire \sr~30_combout ;
wire \sr~31_combout ;
wire \sr~32_combout ;
wire \sr~33_combout ;
wire \sr~34_combout ;
wire \sr~35_combout ;
wire \sr~36_combout ;
wire \sr~37_combout ;
wire \sr~38_combout ;
wire \sr~39_combout ;
wire \sr~40_combout ;
wire \sr~41_combout ;
wire \sr~42_combout ;
wire \sr~43_combout ;
wire \sr~45_combout ;
wire \sr~46_combout ;
wire \sr~47_combout ;
wire \sr~48_combout ;
wire \sr~49_combout ;
wire \sr~50_combout ;
wire \sr~51_combout ;
wire \sr~52_combout ;
wire \sr~53_combout ;
wire \sr~54_combout ;
wire \sr~55_combout ;
wire \sr~56_combout ;
wire \sr~57_combout ;
wire \sr~58_combout ;
wire \sr~59_combout ;
wire \sr~60_combout ;
wire \sr~61_combout ;
wire \sr~62_combout ;
wire \sr~63_combout ;
wire \sr~64_combout ;
wire \sr~65_combout ;
wire \sr~66_combout ;
wire \sr~67_combout ;
wire \sr~68_combout ;
wire \sr~69_combout ;
wire \sr~70_combout ;
wire \sr~73_combout ;
wire \sr~74_combout ;
wire \sr~75_combout ;
wire \sr~76_combout ;
wire \sr~77_combout ;
wire \sr~78_combout ;
wire \sr~79_combout ;
wire \sr~80_combout ;
wire \sr~81_combout ;
wire \sr~82_combout ;


nios_mcu_altera_std_synchronizer_3 the_altera_std_synchronizer2(
	.dreg_0(\the_altera_std_synchronizer2|dreg[0]~q ),
	.din(monitor_ready),
	.clk(altera_internal_jtag));

nios_mcu_altera_std_synchronizer_2 the_altera_std_synchronizer1(
	.dreg_0(\the_altera_std_synchronizer1|dreg[0]~q ),
	.din(hbreak_enabled),
	.clk(altera_internal_jtag));

dffeas \sr[0] (
	.clk(altera_internal_jtag),
	.d(\sr[0]~5_combout ),
	.asdata(\sr~10_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!virtual_state_sdr),
	.ena(vcc),
	.q(sr_0),
	.prn(vcc));
defparam \sr[0] .is_wysiwyg = "true";
defparam \sr[0] .power_up = "low";

dffeas \sr[35] (
	.clk(altera_internal_jtag),
	.d(\sr[35]~6_combout ),
	.asdata(\sr~25_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!virtual_state_sdr),
	.ena(vcc),
	.q(sr_35),
	.prn(vcc));
defparam \sr[35] .is_wysiwyg = "true";
defparam \sr[35] .power_up = "low";

dffeas \sr[31] (
	.clk(altera_internal_jtag),
	.d(\sr[31]~7_combout ),
	.asdata(sr_32),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(virtual_state_sdr),
	.ena(vcc),
	.q(sr_31),
	.prn(vcc));
defparam \sr[31] .is_wysiwyg = "true";
defparam \sr[31] .power_up = "low";

dffeas \sr[7] (
	.clk(altera_internal_jtag),
	.d(\sr[7]~8_combout ),
	.asdata(sr_8),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(virtual_state_sdr),
	.ena(vcc),
	.q(sr_7),
	.prn(vcc));
defparam \sr[7] .is_wysiwyg = "true";
defparam \sr[7] .power_up = "low";

dffeas \sr[15] (
	.clk(altera_internal_jtag),
	.d(\sr[15]~9_combout ),
	.asdata(\sr~72_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!virtual_state_sdr),
	.ena(vcc),
	.q(sr_15),
	.prn(vcc));
defparam \sr[15] .is_wysiwyg = "true";
defparam \sr[15] .power_up = "low";

dffeas \ir_out[0] (
	.clk(altera_internal_jtag),
	.d(\the_altera_std_synchronizer2|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ir_out_0),
	.prn(vcc));
defparam \ir_out[0] .is_wysiwyg = "true";
defparam \ir_out[0] .power_up = "low";

dffeas \ir_out[1] (
	.clk(altera_internal_jtag),
	.d(\the_altera_std_synchronizer1|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ir_out_1),
	.prn(vcc));
defparam \ir_out[1] .is_wysiwyg = "true";
defparam \ir_out[1] .power_up = "low";

dffeas \sr[1] (
	.clk(altera_internal_jtag),
	.d(\sr~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[14]~13_combout ),
	.q(sr_1),
	.prn(vcc));
defparam \sr[1] .is_wysiwyg = "true";
defparam \sr[1] .power_up = "low";

dffeas \sr[2] (
	.clk(altera_internal_jtag),
	.d(\sr~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[14]~13_combout ),
	.q(sr_2),
	.prn(vcc));
defparam \sr[2] .is_wysiwyg = "true";
defparam \sr[2] .power_up = "low";

dffeas \sr[3] (
	.clk(altera_internal_jtag),
	.d(\sr~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[14]~13_combout ),
	.q(sr_3),
	.prn(vcc));
defparam \sr[3] .is_wysiwyg = "true";
defparam \sr[3] .power_up = "low";

dffeas \sr[4] (
	.clk(altera_internal_jtag),
	.d(\sr~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[14]~13_combout ),
	.q(sr_4),
	.prn(vcc));
defparam \sr[4] .is_wysiwyg = "true";
defparam \sr[4] .power_up = "low";

dffeas \sr[36] (
	.clk(altera_internal_jtag),
	.d(\sr~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[37]~21_combout ),
	.q(sr_36),
	.prn(vcc));
defparam \sr[36] .is_wysiwyg = "true";
defparam \sr[36] .power_up = "low";

dffeas \sr[37] (
	.clk(altera_internal_jtag),
	.d(\sr~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[37]~21_combout ),
	.q(sr_37),
	.prn(vcc));
defparam \sr[37] .is_wysiwyg = "true";
defparam \sr[37] .power_up = "low";

dffeas \sr[17] (
	.clk(altera_internal_jtag),
	.d(\sr~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_17),
	.prn(vcc));
defparam \sr[17] .is_wysiwyg = "true";
defparam \sr[17] .power_up = "low";

dffeas \sr[34] (
	.clk(altera_internal_jtag),
	.d(\sr~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_34),
	.prn(vcc));
defparam \sr[34] .is_wysiwyg = "true";
defparam \sr[34] .power_up = "low";

dffeas \sr[5] (
	.clk(altera_internal_jtag),
	.d(\sr~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[14]~13_combout ),
	.q(sr_5),
	.prn(vcc));
defparam \sr[5] .is_wysiwyg = "true";
defparam \sr[5] .power_up = "low";

dffeas \sr[25] (
	.clk(altera_internal_jtag),
	.d(\sr~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_25),
	.prn(vcc));
defparam \sr[25] .is_wysiwyg = "true";
defparam \sr[25] .power_up = "low";

dffeas \sr[21] (
	.clk(altera_internal_jtag),
	.d(\sr~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_21),
	.prn(vcc));
defparam \sr[21] .is_wysiwyg = "true";
defparam \sr[21] .power_up = "low";

dffeas \sr[20] (
	.clk(altera_internal_jtag),
	.d(\sr~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_20),
	.prn(vcc));
defparam \sr[20] .is_wysiwyg = "true";
defparam \sr[20] .power_up = "low";

dffeas \sr[18] (
	.clk(altera_internal_jtag),
	.d(\sr~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_18),
	.prn(vcc));
defparam \sr[18] .is_wysiwyg = "true";
defparam \sr[18] .power_up = "low";

dffeas \sr[33] (
	.clk(altera_internal_jtag),
	.d(\sr~41_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_33),
	.prn(vcc));
defparam \sr[33] .is_wysiwyg = "true";
defparam \sr[33] .power_up = "low";

dffeas \sr[32] (
	.clk(altera_internal_jtag),
	.d(\sr~43_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_32),
	.prn(vcc));
defparam \sr[32] .is_wysiwyg = "true";
defparam \sr[32] .power_up = "low";

dffeas \sr[30] (
	.clk(altera_internal_jtag),
	.d(\sr~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_30),
	.prn(vcc));
defparam \sr[30] .is_wysiwyg = "true";
defparam \sr[30] .power_up = "low";

dffeas \sr[29] (
	.clk(altera_internal_jtag),
	.d(\sr~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_29),
	.prn(vcc));
defparam \sr[29] .is_wysiwyg = "true";
defparam \sr[29] .power_up = "low";

dffeas \sr[28] (
	.clk(altera_internal_jtag),
	.d(\sr~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_28),
	.prn(vcc));
defparam \sr[28] .is_wysiwyg = "true";
defparam \sr[28] .power_up = "low";

dffeas \sr[27] (
	.clk(altera_internal_jtag),
	.d(\sr~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_27),
	.prn(vcc));
defparam \sr[27] .is_wysiwyg = "true";
defparam \sr[27] .power_up = "low";

dffeas \sr[26] (
	.clk(altera_internal_jtag),
	.d(\sr~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_26),
	.prn(vcc));
defparam \sr[26] .is_wysiwyg = "true";
defparam \sr[26] .power_up = "low";

dffeas \sr[6] (
	.clk(altera_internal_jtag),
	.d(\sr~56_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[14]~13_combout ),
	.q(sr_6),
	.prn(vcc));
defparam \sr[6] .is_wysiwyg = "true";
defparam \sr[6] .power_up = "low";

dffeas \sr[19] (
	.clk(altera_internal_jtag),
	.d(\sr~58_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_19),
	.prn(vcc));
defparam \sr[19] .is_wysiwyg = "true";
defparam \sr[19] .power_up = "low";

dffeas \sr[22] (
	.clk(altera_internal_jtag),
	.d(\sr~60_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_22),
	.prn(vcc));
defparam \sr[22] .is_wysiwyg = "true";
defparam \sr[22] .power_up = "low";

dffeas \sr[23] (
	.clk(altera_internal_jtag),
	.d(\sr~62_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_23),
	.prn(vcc));
defparam \sr[23] .is_wysiwyg = "true";
defparam \sr[23] .power_up = "low";

dffeas \sr[16] (
	.clk(altera_internal_jtag),
	.d(\sr~64_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_16),
	.prn(vcc));
defparam \sr[16] .is_wysiwyg = "true";
defparam \sr[16] .power_up = "low";

dffeas \sr[8] (
	.clk(altera_internal_jtag),
	.d(\sr~66_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[14]~13_combout ),
	.q(sr_8),
	.prn(vcc));
defparam \sr[8] .is_wysiwyg = "true";
defparam \sr[8] .power_up = "low";

dffeas \sr[24] (
	.clk(altera_internal_jtag),
	.d(\sr~68_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[33]~29_combout ),
	.q(sr_24),
	.prn(vcc));
defparam \sr[24] .is_wysiwyg = "true";
defparam \sr[24] .power_up = "low";

dffeas \sr[14] (
	.clk(altera_internal_jtag),
	.d(\sr~70_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[14]~13_combout ),
	.q(sr_14),
	.prn(vcc));
defparam \sr[14] .is_wysiwyg = "true";
defparam \sr[14] .power_up = "low";

dffeas \sr[13] (
	.clk(altera_internal_jtag),
	.d(\sr~74_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[14]~13_combout ),
	.q(sr_13),
	.prn(vcc));
defparam \sr[13] .is_wysiwyg = "true";
defparam \sr[13] .power_up = "low";

dffeas \sr[12] (
	.clk(altera_internal_jtag),
	.d(\sr~76_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[14]~13_combout ),
	.q(sr_12),
	.prn(vcc));
defparam \sr[12] .is_wysiwyg = "true";
defparam \sr[12] .power_up = "low";

dffeas \sr[11] (
	.clk(altera_internal_jtag),
	.d(\sr~78_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[14]~13_combout ),
	.q(sr_11),
	.prn(vcc));
defparam \sr[11] .is_wysiwyg = "true";
defparam \sr[11] .power_up = "low";

dffeas \sr[10] (
	.clk(altera_internal_jtag),
	.d(\sr~80_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[14]~13_combout ),
	.q(sr_10),
	.prn(vcc));
defparam \sr[10] .is_wysiwyg = "true";
defparam \sr[10] .power_up = "low";

dffeas \sr[9] (
	.clk(altera_internal_jtag),
	.d(\sr~82_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[14]~13_combout ),
	.q(sr_9),
	.prn(vcc));
defparam \sr[9] .is_wysiwyg = "true";
defparam \sr[9] .power_up = "low";

dffeas \DRsize.000 (
	.clk(altera_internal_jtag),
	.d(vcc),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(virtual_state_uir),
	.q(\DRsize.000~q ),
	.prn(vcc));
defparam \DRsize.000 .is_wysiwyg = "true";
defparam \DRsize.000 .power_up = "low";

cycloneive_lcell_comb \sr[0]~5 (
	.dataa(altera_internal_jtag1),
	.datab(sr_1),
	.datac(gnd),
	.datad(\DRsize.000~q ),
	.cin(gnd),
	.combout(\sr[0]~5_combout ),
	.cout());
defparam \sr[0]~5 .lut_mask = 16'hAACC;
defparam \sr[0]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux37~0 (
	.dataa(irf_reg_0_2),
	.datab(irf_reg_1_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux37~0_combout ),
	.cout());
defparam \Mux37~0 .lut_mask = 16'h7777;
defparam \Mux37~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~10 (
	.dataa(sr_0),
	.datab(virtual_state_cdr),
	.datac(\the_altera_std_synchronizer2|dreg[0]~q ),
	.datad(\Mux37~0_combout ),
	.cin(gnd),
	.combout(\sr~10_combout ),
	.cout());
defparam \sr~10 .lut_mask = 16'hFFB8;
defparam \sr~10 .sum_lutc_input = "datac";

dffeas \DRsize.100 (
	.clk(altera_internal_jtag),
	.d(\Mux37~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(virtual_state_uir),
	.q(\DRsize.100~q ),
	.prn(vcc));
defparam \DRsize.100 .is_wysiwyg = "true";
defparam \DRsize.100 .power_up = "low";

cycloneive_lcell_comb \sr[35]~6 (
	.dataa(sr_36),
	.datab(altera_internal_jtag1),
	.datac(gnd),
	.datad(\DRsize.100~q ),
	.cin(gnd),
	.combout(\sr[35]~6_combout ),
	.cout());
defparam \sr[35]~6 .lut_mask = 16'hAACC;
defparam \sr[35]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~23 (
	.dataa(sr_35),
	.datab(virtual_state_cdr),
	.datac(irf_reg_0_2),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~23_combout ),
	.cout());
defparam \sr~23 .lut_mask = 16'hFFFE;
defparam \sr~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~24 (
	.dataa(state_3),
	.datab(splitter_nodes_receive_1_3),
	.datac(\the_altera_std_synchronizer1|dreg[0]~q ),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\sr~24_combout ),
	.cout());
defparam \sr~24 .lut_mask = 16'hFEFF;
defparam \sr~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~25 (
	.dataa(\sr~23_combout ),
	.datab(\sr~24_combout ),
	.datac(irf_reg_0_2),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~25_combout ),
	.cout());
defparam \sr~25 .lut_mask = 16'hEFFF;
defparam \sr~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr[31]~44 (
	.dataa(irf_reg_0_2),
	.datab(irf_reg_1_2),
	.datac(break_readreg_30),
	.datad(MonDReg_30),
	.cin(gnd),
	.combout(\sr[31]~44_combout ),
	.cout());
defparam \sr[31]~44 .lut_mask = 16'hFFF6;
defparam \sr[31]~44 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr[31]~7 (
	.dataa(sr_31),
	.datab(virtual_state_cdr),
	.datac(irf_reg_0_2),
	.datad(\sr[31]~44_combout ),
	.cin(gnd),
	.combout(\sr[31]~7_combout ),
	.cout());
defparam \sr[31]~7 .lut_mask = 16'hBF8F;
defparam \sr[31]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux30~0 (
	.dataa(break_readreg_6),
	.datab(MonDReg_6),
	.datac(irf_reg_1_2),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\Mux30~0_combout ),
	.cout());
defparam \Mux30~0 .lut_mask = 16'hACFF;
defparam \Mux30~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr[7]~8 (
	.dataa(\Mux30~0_combout ),
	.datab(sr_7),
	.datac(gnd),
	.datad(virtual_state_cdr),
	.cin(gnd),
	.combout(\sr[7]~8_combout ),
	.cout());
defparam \sr[7]~8 .lut_mask = 16'hAACC;
defparam \sr[7]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr[33]~83 (
	.dataa(irf_reg_0_2),
	.datab(irf_reg_1_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sr[33]~83_combout ),
	.cout());
defparam \sr[33]~83 .lut_mask = 16'hEEEE;
defparam \sr[33]~83 .sum_lutc_input = "datac";

dffeas \DRsize.010 (
	.clk(altera_internal_jtag),
	.d(\sr[33]~83_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(virtual_state_uir),
	.q(\DRsize.010~q ),
	.prn(vcc));
defparam \DRsize.010 .is_wysiwyg = "true";
defparam \DRsize.010 .power_up = "low";

cycloneive_lcell_comb \sr[15]~9 (
	.dataa(sr_16),
	.datab(altera_internal_jtag1),
	.datac(gnd),
	.datad(\DRsize.010~q ),
	.cin(gnd),
	.combout(\sr[15]~9_combout ),
	.cout());
defparam \sr[15]~9 .lut_mask = 16'hAACC;
defparam \sr[15]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~71 (
	.dataa(break_readreg_14),
	.datab(MonDReg_14),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~71_combout ),
	.cout());
defparam \sr~71 .lut_mask = 16'hAACC;
defparam \sr~71 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~72 (
	.dataa(sr_15),
	.datab(virtual_state_cdr),
	.datac(\sr~71_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~72_combout ),
	.cout());
defparam \sr~72 .lut_mask = 16'hB8FF;
defparam \sr~72 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~11 (
	.dataa(break_readreg_0),
	.datab(MonDReg_0),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~11_combout ),
	.cout());
defparam \sr~11 .lut_mask = 16'hAACC;
defparam \sr~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~12 (
	.dataa(sr_2),
	.datab(virtual_state_sdr),
	.datac(\sr~11_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~12_combout ),
	.cout());
defparam \sr~12 .lut_mask = 16'hB8FF;
defparam \sr~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr[14]~13 (
	.dataa(splitter_nodes_receive_1_3),
	.datab(state_3),
	.datac(state_4),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\sr[14]~13_combout ),
	.cout());
defparam \sr[14]~13 .lut_mask = 16'hFEFF;
defparam \sr[14]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~14 (
	.dataa(break_readreg_1),
	.datab(MonDReg_1),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~14_combout ),
	.cout());
defparam \sr~14 .lut_mask = 16'hAACC;
defparam \sr~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~15 (
	.dataa(sr_3),
	.datab(virtual_state_sdr),
	.datac(\sr~14_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~15_combout ),
	.cout());
defparam \sr~15 .lut_mask = 16'hB8FF;
defparam \sr~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~16 (
	.dataa(break_readreg_2),
	.datab(MonDReg_2),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~16_combout ),
	.cout());
defparam \sr~16 .lut_mask = 16'hAACC;
defparam \sr~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~17 (
	.dataa(sr_4),
	.datab(virtual_state_sdr),
	.datac(\sr~16_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~17_combout ),
	.cout());
defparam \sr~17 .lut_mask = 16'hB8FF;
defparam \sr~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~18 (
	.dataa(break_readreg_3),
	.datab(MonDReg_3),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~18_combout ),
	.cout());
defparam \sr~18 .lut_mask = 16'hAACC;
defparam \sr~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~19 (
	.dataa(sr_5),
	.datab(virtual_state_sdr),
	.datac(\sr~18_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~19_combout ),
	.cout());
defparam \sr~19 .lut_mask = 16'hB8FF;
defparam \sr~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~20 (
	.dataa(splitter_nodes_receive_1_3),
	.datab(state_4),
	.datac(sr_37),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\sr~20_combout ),
	.cout());
defparam \sr~20 .lut_mask = 16'hFEFF;
defparam \sr~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr[37]~21 (
	.dataa(virtual_state_cdr),
	.datab(irf_reg_0_2),
	.datac(irf_reg_1_2),
	.datad(virtual_state_sdr),
	.cin(gnd),
	.combout(\sr[37]~21_combout ),
	.cout());
defparam \sr[37]~21 .lut_mask = 16'hFF7D;
defparam \sr[37]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~22 (
	.dataa(altera_internal_jtag1),
	.datab(splitter_nodes_receive_1_3),
	.datac(state_4),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\sr~22_combout ),
	.cout());
defparam \sr~22 .lut_mask = 16'hFEFF;
defparam \sr~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~26 (
	.dataa(break_readreg_16),
	.datab(MonDReg_16),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~26_combout ),
	.cout());
defparam \sr~26 .lut_mask = 16'hAACC;
defparam \sr~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~27 (
	.dataa(virtual_state_sdr),
	.datab(irf_reg_0_2),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~27_combout ),
	.cout());
defparam \sr~27 .lut_mask = 16'hEEFF;
defparam \sr~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~28 (
	.dataa(virtual_state_sdr),
	.datab(sr_18),
	.datac(\sr~26_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~28_combout ),
	.cout());
defparam \sr~28 .lut_mask = 16'hFEFF;
defparam \sr~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr[33]~29 (
	.dataa(virtual_state_cdr),
	.datab(irf_reg_0_2),
	.datac(irf_reg_1_2),
	.datad(virtual_state_sdr),
	.cin(gnd),
	.combout(\sr[33]~29_combout ),
	.cout());
defparam \sr[33]~29 .lut_mask = 16'hFF7F;
defparam \sr[33]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~30 (
	.dataa(sr_35),
	.datab(virtual_state_sdr),
	.datac(monitor_error),
	.datad(\Mux37~0_combout ),
	.cin(gnd),
	.combout(\sr~30_combout ),
	.cout());
defparam \sr~30 .lut_mask = 16'hFFB8;
defparam \sr~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~31 (
	.dataa(break_readreg_4),
	.datab(MonDReg_4),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~31_combout ),
	.cout());
defparam \sr~31 .lut_mask = 16'hAACC;
defparam \sr~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~32 (
	.dataa(sr_6),
	.datab(virtual_state_sdr),
	.datac(\sr~31_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~32_combout ),
	.cout());
defparam \sr~32 .lut_mask = 16'hB8FF;
defparam \sr~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~33 (
	.dataa(break_readreg_24),
	.datab(MonDReg_24),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~33_combout ),
	.cout());
defparam \sr~33 .lut_mask = 16'hAACC;
defparam \sr~33 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~34 (
	.dataa(virtual_state_sdr),
	.datab(sr_26),
	.datac(\sr~33_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~34_combout ),
	.cout());
defparam \sr~34 .lut_mask = 16'hFEFF;
defparam \sr~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~35 (
	.dataa(break_readreg_20),
	.datab(MonDReg_20),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~35_combout ),
	.cout());
defparam \sr~35 .lut_mask = 16'hAACC;
defparam \sr~35 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~36 (
	.dataa(virtual_state_sdr),
	.datab(sr_22),
	.datac(\sr~35_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~36_combout ),
	.cout());
defparam \sr~36 .lut_mask = 16'hFEFF;
defparam \sr~36 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~37 (
	.dataa(break_readreg_19),
	.datab(MonDReg_19),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~37_combout ),
	.cout());
defparam \sr~37 .lut_mask = 16'hAACC;
defparam \sr~37 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~38 (
	.dataa(virtual_state_sdr),
	.datab(sr_21),
	.datac(\sr~37_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~38_combout ),
	.cout());
defparam \sr~38 .lut_mask = 16'hFEFF;
defparam \sr~38 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~39 (
	.dataa(break_readreg_17),
	.datab(MonDReg_17),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~39_combout ),
	.cout());
defparam \sr~39 .lut_mask = 16'hAACC;
defparam \sr~39 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~40 (
	.dataa(virtual_state_sdr),
	.datab(sr_19),
	.datac(\sr~39_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~40_combout ),
	.cout());
defparam \sr~40 .lut_mask = 16'hFEFF;
defparam \sr~40 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~41 (
	.dataa(sr_34),
	.datab(virtual_state_sdr),
	.datac(resetlatch),
	.datad(\Mux37~0_combout ),
	.cin(gnd),
	.combout(\sr~41_combout ),
	.cout());
defparam \sr~41 .lut_mask = 16'hFFB8;
defparam \sr~41 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~42 (
	.dataa(break_readreg_31),
	.datab(MonDReg_31),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~42_combout ),
	.cout());
defparam \sr~42 .lut_mask = 16'hAACC;
defparam \sr~42 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~43 (
	.dataa(virtual_state_sdr),
	.datab(sr_33),
	.datac(\sr~42_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~43_combout ),
	.cout());
defparam \sr~43 .lut_mask = 16'hFEFF;
defparam \sr~43 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~45 (
	.dataa(break_readreg_29),
	.datab(MonDReg_29),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~45_combout ),
	.cout());
defparam \sr~45 .lut_mask = 16'hAACC;
defparam \sr~45 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~46 (
	.dataa(virtual_state_sdr),
	.datab(sr_31),
	.datac(\sr~45_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~46_combout ),
	.cout());
defparam \sr~46 .lut_mask = 16'hFEFF;
defparam \sr~46 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~47 (
	.dataa(break_readreg_28),
	.datab(MonDReg_28),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~47_combout ),
	.cout());
defparam \sr~47 .lut_mask = 16'hAACC;
defparam \sr~47 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~48 (
	.dataa(virtual_state_sdr),
	.datab(sr_30),
	.datac(\sr~47_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~48_combout ),
	.cout());
defparam \sr~48 .lut_mask = 16'hFEFF;
defparam \sr~48 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~49 (
	.dataa(break_readreg_27),
	.datab(MonDReg_27),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~49_combout ),
	.cout());
defparam \sr~49 .lut_mask = 16'hAACC;
defparam \sr~49 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~50 (
	.dataa(virtual_state_sdr),
	.datab(sr_29),
	.datac(\sr~49_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~50_combout ),
	.cout());
defparam \sr~50 .lut_mask = 16'hFEFF;
defparam \sr~50 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~51 (
	.dataa(break_readreg_26),
	.datab(MonDReg_26),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~51_combout ),
	.cout());
defparam \sr~51 .lut_mask = 16'hAACC;
defparam \sr~51 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~52 (
	.dataa(virtual_state_sdr),
	.datab(sr_28),
	.datac(\sr~51_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~52_combout ),
	.cout());
defparam \sr~52 .lut_mask = 16'hFEFF;
defparam \sr~52 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~53 (
	.dataa(break_readreg_25),
	.datab(MonDReg_25),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~53_combout ),
	.cout());
defparam \sr~53 .lut_mask = 16'hAACC;
defparam \sr~53 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~54 (
	.dataa(virtual_state_sdr),
	.datab(sr_27),
	.datac(\sr~53_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~54_combout ),
	.cout());
defparam \sr~54 .lut_mask = 16'hFEFF;
defparam \sr~54 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~55 (
	.dataa(break_readreg_5),
	.datab(MonDReg_5),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~55_combout ),
	.cout());
defparam \sr~55 .lut_mask = 16'hAACC;
defparam \sr~55 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~56 (
	.dataa(sr_7),
	.datab(virtual_state_sdr),
	.datac(\sr~55_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~56_combout ),
	.cout());
defparam \sr~56 .lut_mask = 16'hB8FF;
defparam \sr~56 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~57 (
	.dataa(break_readreg_18),
	.datab(MonDReg_18),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~57_combout ),
	.cout());
defparam \sr~57 .lut_mask = 16'hAACC;
defparam \sr~57 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~58 (
	.dataa(virtual_state_sdr),
	.datab(sr_20),
	.datac(\sr~57_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~58_combout ),
	.cout());
defparam \sr~58 .lut_mask = 16'hFEFF;
defparam \sr~58 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~59 (
	.dataa(break_readreg_21),
	.datab(MonDReg_21),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~59_combout ),
	.cout());
defparam \sr~59 .lut_mask = 16'hAACC;
defparam \sr~59 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~60 (
	.dataa(virtual_state_sdr),
	.datab(sr_23),
	.datac(\sr~59_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~60_combout ),
	.cout());
defparam \sr~60 .lut_mask = 16'hFEFF;
defparam \sr~60 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~61 (
	.dataa(break_readreg_22),
	.datab(MonDReg_22),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~61_combout ),
	.cout());
defparam \sr~61 .lut_mask = 16'hAACC;
defparam \sr~61 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~62 (
	.dataa(virtual_state_sdr),
	.datab(sr_24),
	.datac(\sr~61_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~62_combout ),
	.cout());
defparam \sr~62 .lut_mask = 16'hFEFF;
defparam \sr~62 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~63 (
	.dataa(break_readreg_15),
	.datab(MonDReg_15),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~63_combout ),
	.cout());
defparam \sr~63 .lut_mask = 16'hAACC;
defparam \sr~63 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~64 (
	.dataa(virtual_state_sdr),
	.datab(sr_17),
	.datac(\sr~63_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~64_combout ),
	.cout());
defparam \sr~64 .lut_mask = 16'hFEFF;
defparam \sr~64 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~65 (
	.dataa(break_readreg_7),
	.datab(MonDReg_7),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~65_combout ),
	.cout());
defparam \sr~65 .lut_mask = 16'hAACC;
defparam \sr~65 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~66 (
	.dataa(sr_9),
	.datab(virtual_state_sdr),
	.datac(\sr~65_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~66_combout ),
	.cout());
defparam \sr~66 .lut_mask = 16'hB8FF;
defparam \sr~66 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~67 (
	.dataa(break_readreg_23),
	.datab(MonDReg_23),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~67_combout ),
	.cout());
defparam \sr~67 .lut_mask = 16'hAACC;
defparam \sr~67 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~68 (
	.dataa(virtual_state_sdr),
	.datab(sr_25),
	.datac(\sr~67_combout ),
	.datad(\sr~27_combout ),
	.cin(gnd),
	.combout(\sr~68_combout ),
	.cout());
defparam \sr~68 .lut_mask = 16'hFEFF;
defparam \sr~68 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~69 (
	.dataa(break_readreg_13),
	.datab(MonDReg_13),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~69_combout ),
	.cout());
defparam \sr~69 .lut_mask = 16'hAACC;
defparam \sr~69 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~70 (
	.dataa(sr_15),
	.datab(virtual_state_sdr),
	.datac(\sr~69_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~70_combout ),
	.cout());
defparam \sr~70 .lut_mask = 16'hB8FF;
defparam \sr~70 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~73 (
	.dataa(break_readreg_12),
	.datab(MonDReg_12),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~73_combout ),
	.cout());
defparam \sr~73 .lut_mask = 16'hAACC;
defparam \sr~73 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~74 (
	.dataa(sr_14),
	.datab(virtual_state_sdr),
	.datac(\sr~73_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~74_combout ),
	.cout());
defparam \sr~74 .lut_mask = 16'hB8FF;
defparam \sr~74 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~75 (
	.dataa(break_readreg_11),
	.datab(MonDReg_11),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~75_combout ),
	.cout());
defparam \sr~75 .lut_mask = 16'hAACC;
defparam \sr~75 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~76 (
	.dataa(sr_13),
	.datab(virtual_state_sdr),
	.datac(\sr~75_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~76_combout ),
	.cout());
defparam \sr~76 .lut_mask = 16'hB8FF;
defparam \sr~76 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~77 (
	.dataa(break_readreg_10),
	.datab(MonDReg_10),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~77_combout ),
	.cout());
defparam \sr~77 .lut_mask = 16'hAACC;
defparam \sr~77 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~78 (
	.dataa(sr_12),
	.datab(virtual_state_sdr),
	.datac(\sr~77_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~78_combout ),
	.cout());
defparam \sr~78 .lut_mask = 16'hB8FF;
defparam \sr~78 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~79 (
	.dataa(break_readreg_9),
	.datab(MonDReg_9),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~79_combout ),
	.cout());
defparam \sr~79 .lut_mask = 16'hAACC;
defparam \sr~79 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~80 (
	.dataa(sr_11),
	.datab(virtual_state_sdr),
	.datac(\sr~79_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~80_combout ),
	.cout());
defparam \sr~80 .lut_mask = 16'hB8FF;
defparam \sr~80 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~81 (
	.dataa(break_readreg_8),
	.datab(MonDReg_8),
	.datac(gnd),
	.datad(irf_reg_1_2),
	.cin(gnd),
	.combout(\sr~81_combout ),
	.cout());
defparam \sr~81 .lut_mask = 16'hAACC;
defparam \sr~81 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sr~82 (
	.dataa(sr_10),
	.datab(virtual_state_sdr),
	.datac(\sr~81_combout ),
	.datad(irf_reg_0_2),
	.cin(gnd),
	.combout(\sr~82_combout ),
	.cout());
defparam \sr~82 .lut_mask = 16'hB8FF;
defparam \sr~82 .sum_lutc_input = "datac";

endmodule

module nios_mcu_altera_std_synchronizer_2 (
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module nios_mcu_altera_std_synchronizer_3 (
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module nios_mcu_sld_virtual_jtag_basic_1 (
	virtual_state_cdr1,
	virtual_state_sdr,
	virtual_state_uir,
	virtual_state_udr,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3)/* synthesis synthesis_greybox=1 */;
output 	virtual_state_cdr1;
output 	virtual_state_sdr;
output 	virtual_state_uir;
output 	virtual_state_udr;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb virtual_state_cdr(
	.dataa(virtual_ir_scan_reg),
	.datab(gnd),
	.datac(state_3),
	.datad(splitter_nodes_receive_1_3),
	.cin(gnd),
	.combout(virtual_state_cdr1),
	.cout());
defparam virtual_state_cdr.lut_mask = 16'hAFFF;
defparam virtual_state_cdr.sum_lutc_input = "datac";

cycloneive_lcell_comb \virtual_state_sdr~0 (
	.dataa(splitter_nodes_receive_1_3),
	.datab(state_4),
	.datac(gnd),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(virtual_state_sdr),
	.cout());
defparam \virtual_state_sdr~0 .lut_mask = 16'hEEFF;
defparam \virtual_state_sdr~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \virtual_state_uir~0 (
	.dataa(virtual_ir_scan_reg),
	.datab(splitter_nodes_receive_1_3),
	.datac(state_8),
	.datad(gnd),
	.cin(gnd),
	.combout(virtual_state_uir),
	.cout());
defparam \virtual_state_uir~0 .lut_mask = 16'hFEFE;
defparam \virtual_state_uir~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \virtual_state_udr~0 (
	.dataa(splitter_nodes_receive_1_3),
	.datab(state_8),
	.datac(gnd),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(virtual_state_udr),
	.cout());
defparam \virtual_state_udr~0 .lut_mask = 16'hEEFF;
defparam \virtual_state_udr~0 .sum_lutc_input = "datac";

endmodule

module nios_mcu_nios_mcu_nios_cpu_cpu_nios2_avalon_reg (
	r_sync_rst,
	write,
	address_8,
	debugaccess,
	writedata_0,
	address_0,
	address_1,
	address_2,
	address_3,
	address_4,
	address_5,
	address_6,
	address_7,
	Equal0,
	take_action_ocireg,
	oci_ienable_0,
	oci_single_step_mode1,
	monitor_error,
	Equal1,
	oci_reg_readdata_0,
	writedata_3,
	oci_ienable_16,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	write;
input 	address_8;
input 	debugaccess;
input 	writedata_0;
input 	address_0;
input 	address_1;
input 	address_2;
input 	address_3;
input 	address_4;
input 	address_5;
input 	address_6;
input 	address_7;
output 	Equal0;
output 	take_action_ocireg;
output 	oci_ienable_0;
output 	oci_single_step_mode1;
input 	monitor_error;
output 	Equal1;
output 	oci_reg_readdata_0;
input 	writedata_3;
output 	oci_ienable_16;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Equal0~0_combout ;
wire \Equal0~1_combout ;
wire \oci_ienable[0]~0_combout ;
wire \take_action_oci_intr_mask_reg~0_combout ;
wire \oci_single_step_mode~0_combout ;


cycloneive_lcell_comb \Equal0~2 (
	.dataa(\Equal0~0_combout ),
	.datab(\Equal0~1_combout ),
	.datac(gnd),
	.datad(address_0),
	.cin(gnd),
	.combout(Equal0),
	.cout());
defparam \Equal0~2 .lut_mask = 16'hEEFF;
defparam \Equal0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \take_action_ocireg~0 (
	.dataa(write),
	.datab(debugaccess),
	.datac(Equal0),
	.datad(gnd),
	.cin(gnd),
	.combout(take_action_ocireg),
	.cout());
defparam \take_action_ocireg~0 .lut_mask = 16'hFEFE;
defparam \take_action_ocireg~0 .sum_lutc_input = "datac";

dffeas \oci_ienable[0] (
	.clk(clk_clk),
	.d(\oci_ienable[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_action_oci_intr_mask_reg~0_combout ),
	.q(oci_ienable_0),
	.prn(vcc));
defparam \oci_ienable[0] .is_wysiwyg = "true";
defparam \oci_ienable[0] .power_up = "low";

dffeas oci_single_step_mode(
	.clk(clk_clk),
	.d(\oci_single_step_mode~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(oci_single_step_mode1),
	.prn(vcc));
defparam oci_single_step_mode.is_wysiwyg = "true";
defparam oci_single_step_mode.power_up = "low";

cycloneive_lcell_comb \Equal1~0 (
	.dataa(address_0),
	.datab(\Equal0~0_combout ),
	.datac(\Equal0~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(Equal1),
	.cout());
defparam \Equal1~0 .lut_mask = 16'hFEFE;
defparam \Equal1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \oci_reg_readdata[0]~0 (
	.dataa(monitor_error),
	.datab(Equal0),
	.datac(Equal1),
	.datad(oci_ienable_0),
	.cin(gnd),
	.combout(oci_reg_readdata_0),
	.cout());
defparam \oci_reg_readdata[0]~0 .lut_mask = 16'hB8FF;
defparam \oci_reg_readdata[0]~0 .sum_lutc_input = "datac";

dffeas \oci_ienable[16] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_action_oci_intr_mask_reg~0_combout ),
	.q(oci_ienable_16),
	.prn(vcc));
defparam \oci_ienable[16] .is_wysiwyg = "true";
defparam \oci_ienable[16] .power_up = "low";

cycloneive_lcell_comb \Equal0~0 (
	.dataa(address_8),
	.datab(address_5),
	.datac(address_6),
	.datad(address_7),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hBFFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~1 (
	.dataa(address_1),
	.datab(address_2),
	.datac(address_3),
	.datad(address_4),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'h7FFF;
defparam \Equal0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \oci_ienable[0]~0 (
	.dataa(writedata_0),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\oci_ienable[0]~0_combout ),
	.cout());
defparam \oci_ienable[0]~0 .lut_mask = 16'h5555;
defparam \oci_ienable[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \take_action_oci_intr_mask_reg~0 (
	.dataa(write),
	.datab(debugaccess),
	.datac(Equal1),
	.datad(gnd),
	.cin(gnd),
	.combout(\take_action_oci_intr_mask_reg~0_combout ),
	.cout());
defparam \take_action_oci_intr_mask_reg~0 .lut_mask = 16'hFEFE;
defparam \take_action_oci_intr_mask_reg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \oci_single_step_mode~0 (
	.dataa(writedata_3),
	.datab(oci_single_step_mode1),
	.datac(gnd),
	.datad(take_action_ocireg),
	.cin(gnd),
	.combout(\oci_single_step_mode~0_combout ),
	.cout());
defparam \oci_single_step_mode~0 .lut_mask = 16'hAACC;
defparam \oci_single_step_mode~0 .sum_lutc_input = "datac";

endmodule

module nios_mcu_nios_mcu_nios_cpu_cpu_nios2_oci_break (
	break_readreg_0,
	break_readreg_1,
	jdo_0,
	jdo_36,
	jdo_37,
	ir_0,
	ir_1,
	enable_action_strobe,
	jdo_3,
	jdo_17,
	break_readreg_2,
	jdo_1,
	jdo_4,
	jdo_25,
	jdo_21,
	jdo_20,
	jdo_31,
	jdo_30,
	jdo_29,
	jdo_28,
	jdo_27,
	jdo_26,
	break_readreg_3,
	jdo_2,
	jdo_5,
	jdo_19,
	jdo_18,
	break_readreg_16,
	break_readreg_4,
	jdo_6,
	break_readreg_24,
	break_readreg_20,
	break_readreg_19,
	jdo_23,
	break_readreg_17,
	jdo_16,
	break_readreg_31,
	break_readreg_30,
	break_readreg_29,
	break_readreg_28,
	break_readreg_27,
	break_readreg_26,
	break_readreg_25,
	break_readreg_5,
	jdo_7,
	jdo_24,
	break_readreg_18,
	break_readreg_21,
	jdo_22,
	jdo_14,
	jdo_15,
	jdo_8,
	jdo_13,
	jdo_12,
	jdo_11,
	jdo_10,
	jdo_9,
	break_readreg_6,
	break_readreg_22,
	break_readreg_15,
	break_readreg_7,
	break_readreg_23,
	break_readreg_13,
	break_readreg_14,
	break_readreg_12,
	break_readreg_11,
	break_readreg_10,
	break_readreg_9,
	break_readreg_8,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	break_readreg_0;
output 	break_readreg_1;
input 	jdo_0;
input 	jdo_36;
input 	jdo_37;
input 	ir_0;
input 	ir_1;
input 	enable_action_strobe;
input 	jdo_3;
input 	jdo_17;
output 	break_readreg_2;
input 	jdo_1;
input 	jdo_4;
input 	jdo_25;
input 	jdo_21;
input 	jdo_20;
input 	jdo_31;
input 	jdo_30;
input 	jdo_29;
input 	jdo_28;
input 	jdo_27;
input 	jdo_26;
output 	break_readreg_3;
input 	jdo_2;
input 	jdo_5;
input 	jdo_19;
input 	jdo_18;
output 	break_readreg_16;
output 	break_readreg_4;
input 	jdo_6;
output 	break_readreg_24;
output 	break_readreg_20;
output 	break_readreg_19;
input 	jdo_23;
output 	break_readreg_17;
input 	jdo_16;
output 	break_readreg_31;
output 	break_readreg_30;
output 	break_readreg_29;
output 	break_readreg_28;
output 	break_readreg_27;
output 	break_readreg_26;
output 	break_readreg_25;
output 	break_readreg_5;
input 	jdo_7;
input 	jdo_24;
output 	break_readreg_18;
output 	break_readreg_21;
input 	jdo_22;
input 	jdo_14;
input 	jdo_15;
input 	jdo_8;
input 	jdo_13;
input 	jdo_12;
input 	jdo_11;
input 	jdo_10;
input 	jdo_9;
output 	break_readreg_6;
output 	break_readreg_22;
output 	break_readreg_15;
output 	break_readreg_7;
output 	break_readreg_23;
output 	break_readreg_13;
output 	break_readreg_14;
output 	break_readreg_12;
output 	break_readreg_11;
output 	break_readreg_10;
output 	break_readreg_9;
output 	break_readreg_8;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \break_readreg~0_combout ;
wire \break_readreg[19]~1_combout ;
wire \break_readreg~2_combout ;
wire \break_readreg~3_combout ;
wire \break_readreg~4_combout ;
wire \break_readreg~5_combout ;
wire \break_readreg~6_combout ;
wire \break_readreg~7_combout ;
wire \break_readreg~8_combout ;
wire \break_readreg~9_combout ;
wire \break_readreg~10_combout ;
wire \break_readreg~11_combout ;
wire \break_readreg~12_combout ;
wire \break_readreg~13_combout ;
wire \break_readreg~14_combout ;
wire \break_readreg~15_combout ;
wire \break_readreg~16_combout ;
wire \break_readreg~17_combout ;
wire \break_readreg~18_combout ;
wire \break_readreg~19_combout ;
wire \break_readreg~20_combout ;
wire \break_readreg~21_combout ;
wire \break_readreg~22_combout ;
wire \break_readreg~23_combout ;
wire \break_readreg~24_combout ;
wire \break_readreg~25_combout ;
wire \break_readreg~26_combout ;
wire \break_readreg~27_combout ;
wire \break_readreg~28_combout ;
wire \break_readreg~29_combout ;
wire \break_readreg~30_combout ;
wire \break_readreg~31_combout ;
wire \break_readreg~32_combout ;


dffeas \break_readreg[0] (
	.clk(clk_clk),
	.d(\break_readreg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_0),
	.prn(vcc));
defparam \break_readreg[0] .is_wysiwyg = "true";
defparam \break_readreg[0] .power_up = "low";

dffeas \break_readreg[1] (
	.clk(clk_clk),
	.d(\break_readreg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_1),
	.prn(vcc));
defparam \break_readreg[1] .is_wysiwyg = "true";
defparam \break_readreg[1] .power_up = "low";

dffeas \break_readreg[2] (
	.clk(clk_clk),
	.d(\break_readreg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_2),
	.prn(vcc));
defparam \break_readreg[2] .is_wysiwyg = "true";
defparam \break_readreg[2] .power_up = "low";

dffeas \break_readreg[3] (
	.clk(clk_clk),
	.d(\break_readreg~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_3),
	.prn(vcc));
defparam \break_readreg[3] .is_wysiwyg = "true";
defparam \break_readreg[3] .power_up = "low";

dffeas \break_readreg[16] (
	.clk(clk_clk),
	.d(\break_readreg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_16),
	.prn(vcc));
defparam \break_readreg[16] .is_wysiwyg = "true";
defparam \break_readreg[16] .power_up = "low";

dffeas \break_readreg[4] (
	.clk(clk_clk),
	.d(\break_readreg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_4),
	.prn(vcc));
defparam \break_readreg[4] .is_wysiwyg = "true";
defparam \break_readreg[4] .power_up = "low";

dffeas \break_readreg[24] (
	.clk(clk_clk),
	.d(\break_readreg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_24),
	.prn(vcc));
defparam \break_readreg[24] .is_wysiwyg = "true";
defparam \break_readreg[24] .power_up = "low";

dffeas \break_readreg[20] (
	.clk(clk_clk),
	.d(\break_readreg~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_20),
	.prn(vcc));
defparam \break_readreg[20] .is_wysiwyg = "true";
defparam \break_readreg[20] .power_up = "low";

dffeas \break_readreg[19] (
	.clk(clk_clk),
	.d(\break_readreg~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_19),
	.prn(vcc));
defparam \break_readreg[19] .is_wysiwyg = "true";
defparam \break_readreg[19] .power_up = "low";

dffeas \break_readreg[17] (
	.clk(clk_clk),
	.d(\break_readreg~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_17),
	.prn(vcc));
defparam \break_readreg[17] .is_wysiwyg = "true";
defparam \break_readreg[17] .power_up = "low";

dffeas \break_readreg[31] (
	.clk(clk_clk),
	.d(\break_readreg~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_31),
	.prn(vcc));
defparam \break_readreg[31] .is_wysiwyg = "true";
defparam \break_readreg[31] .power_up = "low";

dffeas \break_readreg[30] (
	.clk(clk_clk),
	.d(\break_readreg~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_30),
	.prn(vcc));
defparam \break_readreg[30] .is_wysiwyg = "true";
defparam \break_readreg[30] .power_up = "low";

dffeas \break_readreg[29] (
	.clk(clk_clk),
	.d(\break_readreg~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_29),
	.prn(vcc));
defparam \break_readreg[29] .is_wysiwyg = "true";
defparam \break_readreg[29] .power_up = "low";

dffeas \break_readreg[28] (
	.clk(clk_clk),
	.d(\break_readreg~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_28),
	.prn(vcc));
defparam \break_readreg[28] .is_wysiwyg = "true";
defparam \break_readreg[28] .power_up = "low";

dffeas \break_readreg[27] (
	.clk(clk_clk),
	.d(\break_readreg~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_27),
	.prn(vcc));
defparam \break_readreg[27] .is_wysiwyg = "true";
defparam \break_readreg[27] .power_up = "low";

dffeas \break_readreg[26] (
	.clk(clk_clk),
	.d(\break_readreg~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_26),
	.prn(vcc));
defparam \break_readreg[26] .is_wysiwyg = "true";
defparam \break_readreg[26] .power_up = "low";

dffeas \break_readreg[25] (
	.clk(clk_clk),
	.d(\break_readreg~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_25),
	.prn(vcc));
defparam \break_readreg[25] .is_wysiwyg = "true";
defparam \break_readreg[25] .power_up = "low";

dffeas \break_readreg[5] (
	.clk(clk_clk),
	.d(\break_readreg~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_5),
	.prn(vcc));
defparam \break_readreg[5] .is_wysiwyg = "true";
defparam \break_readreg[5] .power_up = "low";

dffeas \break_readreg[18] (
	.clk(clk_clk),
	.d(\break_readreg~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_18),
	.prn(vcc));
defparam \break_readreg[18] .is_wysiwyg = "true";
defparam \break_readreg[18] .power_up = "low";

dffeas \break_readreg[21] (
	.clk(clk_clk),
	.d(\break_readreg~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_21),
	.prn(vcc));
defparam \break_readreg[21] .is_wysiwyg = "true";
defparam \break_readreg[21] .power_up = "low";

dffeas \break_readreg[6] (
	.clk(clk_clk),
	.d(\break_readreg~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_6),
	.prn(vcc));
defparam \break_readreg[6] .is_wysiwyg = "true";
defparam \break_readreg[6] .power_up = "low";

dffeas \break_readreg[22] (
	.clk(clk_clk),
	.d(\break_readreg~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_22),
	.prn(vcc));
defparam \break_readreg[22] .is_wysiwyg = "true";
defparam \break_readreg[22] .power_up = "low";

dffeas \break_readreg[15] (
	.clk(clk_clk),
	.d(\break_readreg~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_15),
	.prn(vcc));
defparam \break_readreg[15] .is_wysiwyg = "true";
defparam \break_readreg[15] .power_up = "low";

dffeas \break_readreg[7] (
	.clk(clk_clk),
	.d(\break_readreg~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_7),
	.prn(vcc));
defparam \break_readreg[7] .is_wysiwyg = "true";
defparam \break_readreg[7] .power_up = "low";

dffeas \break_readreg[23] (
	.clk(clk_clk),
	.d(\break_readreg~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_23),
	.prn(vcc));
defparam \break_readreg[23] .is_wysiwyg = "true";
defparam \break_readreg[23] .power_up = "low";

dffeas \break_readreg[13] (
	.clk(clk_clk),
	.d(\break_readreg~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_13),
	.prn(vcc));
defparam \break_readreg[13] .is_wysiwyg = "true";
defparam \break_readreg[13] .power_up = "low";

dffeas \break_readreg[14] (
	.clk(clk_clk),
	.d(\break_readreg~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_14),
	.prn(vcc));
defparam \break_readreg[14] .is_wysiwyg = "true";
defparam \break_readreg[14] .power_up = "low";

dffeas \break_readreg[12] (
	.clk(clk_clk),
	.d(\break_readreg~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_12),
	.prn(vcc));
defparam \break_readreg[12] .is_wysiwyg = "true";
defparam \break_readreg[12] .power_up = "low";

dffeas \break_readreg[11] (
	.clk(clk_clk),
	.d(\break_readreg~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_11),
	.prn(vcc));
defparam \break_readreg[11] .is_wysiwyg = "true";
defparam \break_readreg[11] .power_up = "low";

dffeas \break_readreg[10] (
	.clk(clk_clk),
	.d(\break_readreg~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_10),
	.prn(vcc));
defparam \break_readreg[10] .is_wysiwyg = "true";
defparam \break_readreg[10] .power_up = "low";

dffeas \break_readreg[9] (
	.clk(clk_clk),
	.d(\break_readreg~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_9),
	.prn(vcc));
defparam \break_readreg[9] .is_wysiwyg = "true";
defparam \break_readreg[9] .power_up = "low";

dffeas \break_readreg[8] (
	.clk(clk_clk),
	.d(\break_readreg~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\break_readreg[19]~1_combout ),
	.q(break_readreg_8),
	.prn(vcc));
defparam \break_readreg[8] .is_wysiwyg = "true";
defparam \break_readreg[8] .power_up = "low";

cycloneive_lcell_comb \break_readreg~0 (
	.dataa(jdo_0),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(gnd),
	.cin(gnd),
	.combout(\break_readreg~0_combout ),
	.cout());
defparam \break_readreg~0 .lut_mask = 16'hFEFE;
defparam \break_readreg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg[19]~1 (
	.dataa(ir_0),
	.datab(gnd),
	.datac(ir_1),
	.datad(enable_action_strobe),
	.cin(gnd),
	.combout(\break_readreg[19]~1_combout ),
	.cout());
defparam \break_readreg[19]~1 .lut_mask = 16'hFFF5;
defparam \break_readreg[19]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~2 (
	.dataa(jdo_1),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(gnd),
	.cin(gnd),
	.combout(\break_readreg~2_combout ),
	.cout());
defparam \break_readreg~2 .lut_mask = 16'hFEFE;
defparam \break_readreg~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~3 (
	.dataa(jdo_2),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(gnd),
	.cin(gnd),
	.combout(\break_readreg~3_combout ),
	.cout());
defparam \break_readreg~3 .lut_mask = 16'hFEFE;
defparam \break_readreg~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~4 (
	.dataa(jdo_3),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~4_combout ),
	.cout());
defparam \break_readreg~4 .lut_mask = 16'hFEFF;
defparam \break_readreg~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~5 (
	.dataa(jdo_16),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~5_combout ),
	.cout());
defparam \break_readreg~5 .lut_mask = 16'hFEFF;
defparam \break_readreg~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~6 (
	.dataa(jdo_4),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~6_combout ),
	.cout());
defparam \break_readreg~6 .lut_mask = 16'hFEFF;
defparam \break_readreg~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~7 (
	.dataa(jdo_24),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~7_combout ),
	.cout());
defparam \break_readreg~7 .lut_mask = 16'hFEFF;
defparam \break_readreg~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~8 (
	.dataa(jdo_20),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~8_combout ),
	.cout());
defparam \break_readreg~8 .lut_mask = 16'hFEFF;
defparam \break_readreg~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~9 (
	.dataa(jdo_19),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~9_combout ),
	.cout());
defparam \break_readreg~9 .lut_mask = 16'hFEFF;
defparam \break_readreg~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~10 (
	.dataa(jdo_17),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~10_combout ),
	.cout());
defparam \break_readreg~10 .lut_mask = 16'hFEFF;
defparam \break_readreg~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~11 (
	.dataa(jdo_31),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~11_combout ),
	.cout());
defparam \break_readreg~11 .lut_mask = 16'hFEFF;
defparam \break_readreg~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~12 (
	.dataa(jdo_30),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~12_combout ),
	.cout());
defparam \break_readreg~12 .lut_mask = 16'hFEFF;
defparam \break_readreg~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~13 (
	.dataa(jdo_29),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~13_combout ),
	.cout());
defparam \break_readreg~13 .lut_mask = 16'hFEFF;
defparam \break_readreg~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~14 (
	.dataa(jdo_28),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~14_combout ),
	.cout());
defparam \break_readreg~14 .lut_mask = 16'hFEFF;
defparam \break_readreg~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~15 (
	.dataa(jdo_27),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~15_combout ),
	.cout());
defparam \break_readreg~15 .lut_mask = 16'hFEFF;
defparam \break_readreg~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~16 (
	.dataa(jdo_26),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~16_combout ),
	.cout());
defparam \break_readreg~16 .lut_mask = 16'hFEFF;
defparam \break_readreg~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~17 (
	.dataa(jdo_25),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~17_combout ),
	.cout());
defparam \break_readreg~17 .lut_mask = 16'hFEFF;
defparam \break_readreg~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~18 (
	.dataa(jdo_5),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~18_combout ),
	.cout());
defparam \break_readreg~18 .lut_mask = 16'hFEFF;
defparam \break_readreg~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~19 (
	.dataa(jdo_18),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~19_combout ),
	.cout());
defparam \break_readreg~19 .lut_mask = 16'hFEFF;
defparam \break_readreg~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~20 (
	.dataa(jdo_21),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~20_combout ),
	.cout());
defparam \break_readreg~20 .lut_mask = 16'hFEFF;
defparam \break_readreg~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~21 (
	.dataa(jdo_6),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~21_combout ),
	.cout());
defparam \break_readreg~21 .lut_mask = 16'hFEFF;
defparam \break_readreg~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~22 (
	.dataa(jdo_22),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~22_combout ),
	.cout());
defparam \break_readreg~22 .lut_mask = 16'hFEFF;
defparam \break_readreg~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~23 (
	.dataa(jdo_15),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~23_combout ),
	.cout());
defparam \break_readreg~23 .lut_mask = 16'hFEFF;
defparam \break_readreg~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~24 (
	.dataa(jdo_7),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~24_combout ),
	.cout());
defparam \break_readreg~24 .lut_mask = 16'hFEFF;
defparam \break_readreg~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~25 (
	.dataa(jdo_23),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~25_combout ),
	.cout());
defparam \break_readreg~25 .lut_mask = 16'hFEFF;
defparam \break_readreg~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~26 (
	.dataa(jdo_13),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~26_combout ),
	.cout());
defparam \break_readreg~26 .lut_mask = 16'hFEFF;
defparam \break_readreg~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~27 (
	.dataa(jdo_14),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~27_combout ),
	.cout());
defparam \break_readreg~27 .lut_mask = 16'hFEFF;
defparam \break_readreg~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~28 (
	.dataa(jdo_12),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~28_combout ),
	.cout());
defparam \break_readreg~28 .lut_mask = 16'hFEFF;
defparam \break_readreg~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~29 (
	.dataa(jdo_11),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~29_combout ),
	.cout());
defparam \break_readreg~29 .lut_mask = 16'hFEFF;
defparam \break_readreg~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~30 (
	.dataa(jdo_10),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~30_combout ),
	.cout());
defparam \break_readreg~30 .lut_mask = 16'hFEFF;
defparam \break_readreg~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~31 (
	.dataa(jdo_9),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~31_combout ),
	.cout());
defparam \break_readreg~31 .lut_mask = 16'hFEFF;
defparam \break_readreg~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \break_readreg~32 (
	.dataa(jdo_8),
	.datab(jdo_36),
	.datac(jdo_37),
	.datad(\break_readreg[19]~1_combout ),
	.cin(gnd),
	.combout(\break_readreg~32_combout ),
	.cout());
defparam \break_readreg~32 .lut_mask = 16'hFEFF;
defparam \break_readreg~32 .sum_lutc_input = "datac";

endmodule

module nios_mcu_nios_mcu_nios_cpu_cpu_nios2_oci_debug (
	jtag_break1,
	r_sync_rst,
	monitor_ready1,
	take_action_ocimem_a,
	jdo_34,
	writedata_0,
	take_action_ocireg,
	jdo_25,
	jdo_21,
	jdo_20,
	take_action_ocimem_a1,
	writedata_1,
	monitor_error1,
	jdo_19,
	jdo_18,
	monitor_go1,
	jdo_23,
	resetlatch1,
	jdo_24,
	state_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	jtag_break1;
input 	r_sync_rst;
output 	monitor_ready1;
input 	take_action_ocimem_a;
input 	jdo_34;
input 	writedata_0;
input 	take_action_ocireg;
input 	jdo_25;
input 	jdo_21;
input 	jdo_20;
input 	take_action_ocimem_a1;
input 	writedata_1;
output 	monitor_error1;
input 	jdo_19;
input 	jdo_18;
output 	monitor_go1;
input 	jdo_23;
output 	resetlatch1;
input 	jdo_24;
input 	state_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_altera_std_synchronizer|dreg[0]~q ;
wire \break_on_reset~0_combout ;
wire \break_on_reset~q ;
wire \jtag_break~0_combout ;
wire \jtag_break~1_combout ;
wire \always1~0_combout ;
wire \monitor_ready~0_combout ;
wire \monitor_error~0_combout ;
wire \monitor_go~0_combout ;
wire \resetlatch~0_combout ;


nios_mcu_altera_std_synchronizer_4 the_altera_std_synchronizer(
	.din(r_sync_rst),
	.dreg_0(\the_altera_std_synchronizer|dreg[0]~q ),
	.clk(clk_clk));

dffeas jtag_break(
	.clk(clk_clk),
	.d(\jtag_break~0_combout ),
	.asdata(\jtag_break~1_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a1),
	.ena(vcc),
	.q(jtag_break1),
	.prn(vcc));
defparam jtag_break.is_wysiwyg = "true";
defparam jtag_break.power_up = "low";

dffeas monitor_ready(
	.clk(clk_clk),
	.d(\monitor_ready~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(monitor_ready1),
	.prn(vcc));
defparam monitor_ready.is_wysiwyg = "true";
defparam monitor_ready.power_up = "low";

dffeas monitor_error(
	.clk(clk_clk),
	.d(\monitor_error~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(monitor_error1),
	.prn(vcc));
defparam monitor_error.is_wysiwyg = "true";
defparam monitor_error.power_up = "low";

dffeas monitor_go(
	.clk(clk_clk),
	.d(\monitor_go~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(monitor_go1),
	.prn(vcc));
defparam monitor_go.is_wysiwyg = "true";
defparam monitor_go.power_up = "low";

dffeas resetlatch(
	.clk(clk_clk),
	.d(\resetlatch~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(resetlatch1),
	.prn(vcc));
defparam resetlatch.is_wysiwyg = "true";
defparam resetlatch.power_up = "low";

cycloneive_lcell_comb \break_on_reset~0 (
	.dataa(jdo_19),
	.datab(\break_on_reset~q ),
	.datac(take_action_ocimem_a1),
	.datad(jdo_18),
	.cin(gnd),
	.combout(\break_on_reset~0_combout ),
	.cout());
defparam \break_on_reset~0 .lut_mask = 16'hACFF;
defparam \break_on_reset~0 .sum_lutc_input = "datac";

dffeas break_on_reset(
	.clk(clk_clk),
	.d(\break_on_reset~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\break_on_reset~q ),
	.prn(vcc));
defparam break_on_reset.is_wysiwyg = "true";
defparam break_on_reset.power_up = "low";

cycloneive_lcell_comb \jtag_break~0 (
	.dataa(jtag_break1),
	.datab(\break_on_reset~q ),
	.datac(gnd),
	.datad(\the_altera_std_synchronizer|dreg[0]~q ),
	.cin(gnd),
	.combout(\jtag_break~0_combout ),
	.cout());
defparam \jtag_break~0 .lut_mask = 16'hAACC;
defparam \jtag_break~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \jtag_break~1 (
	.dataa(jdo_21),
	.datab(jtag_break1),
	.datac(gnd),
	.datad(jdo_20),
	.cin(gnd),
	.combout(\jtag_break~1_combout ),
	.cout());
defparam \jtag_break~1 .lut_mask = 16'hEEFF;
defparam \jtag_break~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always1~0 (
	.dataa(take_action_ocimem_a),
	.datab(jdo_34),
	.datac(jdo_25),
	.datad(gnd),
	.cin(gnd),
	.combout(\always1~0_combout ),
	.cout());
defparam \always1~0 .lut_mask = 16'hFEFE;
defparam \always1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \monitor_ready~0 (
	.dataa(monitor_ready1),
	.datab(writedata_0),
	.datac(take_action_ocireg),
	.datad(\always1~0_combout ),
	.cin(gnd),
	.combout(\monitor_ready~0_combout ),
	.cout());
defparam \monitor_ready~0 .lut_mask = 16'hFEFF;
defparam \monitor_ready~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \monitor_error~0 (
	.dataa(monitor_error1),
	.datab(take_action_ocireg),
	.datac(writedata_1),
	.datad(\always1~0_combout ),
	.cin(gnd),
	.combout(\monitor_error~0_combout ),
	.cout());
defparam \monitor_error~0 .lut_mask = 16'hFEFF;
defparam \monitor_error~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \monitor_go~0 (
	.dataa(take_action_ocimem_a1),
	.datab(jdo_23),
	.datac(monitor_go1),
	.datad(state_1),
	.cin(gnd),
	.combout(\monitor_go~0_combout ),
	.cout());
defparam \monitor_go~0 .lut_mask = 16'hFEFF;
defparam \monitor_go~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \resetlatch~0 (
	.dataa(resetlatch1),
	.datab(\the_altera_std_synchronizer|dreg[0]~q ),
	.datac(jdo_24),
	.datad(take_action_ocimem_a1),
	.cin(gnd),
	.combout(\resetlatch~0_combout ),
	.cout());
defparam \resetlatch~0 .lut_mask = 16'hEFFF;
defparam \resetlatch~0 .sum_lutc_input = "datac";

endmodule

module nios_mcu_altera_std_synchronizer_4 (
	din,
	dreg_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	din;
output 	dreg_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module nios_mcu_nios_mcu_nios_cpu_cpu_nios2_ocimem (
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_22,
	q_a_23,
	q_a_24,
	q_a_25,
	q_a_26,
	q_a_11,
	q_a_13,
	q_a_16,
	q_a_12,
	q_a_3,
	q_a_5,
	q_a_4,
	q_a_14,
	q_a_15,
	q_a_18,
	q_a_17,
	q_a_10,
	q_a_9,
	q_a_8,
	q_a_7,
	q_a_6,
	q_a_21,
	q_a_19,
	q_a_20,
	MonDReg_4,
	MonDReg_12,
	MonDReg_5,
	MonDReg_18,
	q_a_27,
	q_a_28,
	q_a_29,
	q_a_30,
	q_a_31,
	MonDReg_8,
	MonDReg_29,
	waitrequest1,
	MonDReg_0,
	write,
	address_8,
	read,
	MonDReg_1,
	jdo_3,
	jdo_35,
	take_action_ocimem_b,
	take_action_ocimem_a,
	jdo_17,
	take_action_ocimem_a1,
	jdo_34,
	MonDReg_2,
	jdo_4,
	debugaccess,
	r_early_rst,
	writedata_0,
	address_0,
	address_1,
	address_2,
	address_3,
	address_4,
	address_5,
	address_6,
	address_7,
	byteenable_0,
	jdo_25,
	jdo_21,
	jdo_20,
	jdo_33,
	jdo_32,
	jdo_31,
	jdo_30,
	jdo_29,
	jdo_28,
	jdo_27,
	jdo_26,
	MonDReg_3,
	jdo_5,
	writedata_1,
	jdo_19,
	jdo_18,
	writedata_3,
	MonDReg_16,
	jdo_6,
	writedata_2,
	MonDReg_24,
	MonDReg_20,
	MonDReg_19,
	MonDReg_22,
	writedata_22,
	byteenable_2,
	MonDReg_23,
	writedata_23,
	writedata_24,
	byteenable_3,
	MonDReg_25,
	writedata_25,
	MonDReg_26,
	writedata_26,
	MonDReg_11,
	writedata_11,
	byteenable_1,
	MonDReg_13,
	writedata_13,
	writedata_16,
	writedata_12,
	jdo_23,
	writedata_5,
	writedata_4,
	MonDReg_14,
	writedata_14,
	MonDReg_15,
	writedata_15,
	writedata_18,
	MonDReg_17,
	writedata_17,
	MonDReg_10,
	writedata_10,
	MonDReg_9,
	writedata_9,
	writedata_8,
	MonDReg_7,
	writedata_7,
	MonDReg_6,
	writedata_6,
	MonDReg_21,
	writedata_21,
	writedata_19,
	writedata_20,
	jdo_16,
	MonDReg_31,
	MonDReg_30,
	MonDReg_28,
	MonDReg_27,
	jdo_7,
	jdo_24,
	jdo_22,
	jdo_14,
	jdo_15,
	jdo_8,
	writedata_27,
	writedata_28,
	writedata_29,
	writedata_30,
	writedata_31,
	jdo_13,
	jdo_12,
	jdo_11,
	jdo_10,
	jdo_9,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_22;
output 	q_a_23;
output 	q_a_24;
output 	q_a_25;
output 	q_a_26;
output 	q_a_11;
output 	q_a_13;
output 	q_a_16;
output 	q_a_12;
output 	q_a_3;
output 	q_a_5;
output 	q_a_4;
output 	q_a_14;
output 	q_a_15;
output 	q_a_18;
output 	q_a_17;
output 	q_a_10;
output 	q_a_9;
output 	q_a_8;
output 	q_a_7;
output 	q_a_6;
output 	q_a_21;
output 	q_a_19;
output 	q_a_20;
output 	MonDReg_4;
output 	MonDReg_12;
output 	MonDReg_5;
output 	MonDReg_18;
output 	q_a_27;
output 	q_a_28;
output 	q_a_29;
output 	q_a_30;
output 	q_a_31;
output 	MonDReg_8;
output 	MonDReg_29;
output 	waitrequest1;
output 	MonDReg_0;
input 	write;
input 	address_8;
input 	read;
output 	MonDReg_1;
input 	jdo_3;
input 	jdo_35;
input 	take_action_ocimem_b;
input 	take_action_ocimem_a;
input 	jdo_17;
input 	take_action_ocimem_a1;
input 	jdo_34;
output 	MonDReg_2;
input 	jdo_4;
input 	debugaccess;
input 	r_early_rst;
input 	writedata_0;
input 	address_0;
input 	address_1;
input 	address_2;
input 	address_3;
input 	address_4;
input 	address_5;
input 	address_6;
input 	address_7;
input 	byteenable_0;
input 	jdo_25;
input 	jdo_21;
input 	jdo_20;
input 	jdo_33;
input 	jdo_32;
input 	jdo_31;
input 	jdo_30;
input 	jdo_29;
input 	jdo_28;
input 	jdo_27;
input 	jdo_26;
output 	MonDReg_3;
input 	jdo_5;
input 	writedata_1;
input 	jdo_19;
input 	jdo_18;
input 	writedata_3;
output 	MonDReg_16;
input 	jdo_6;
input 	writedata_2;
output 	MonDReg_24;
output 	MonDReg_20;
output 	MonDReg_19;
output 	MonDReg_22;
input 	writedata_22;
input 	byteenable_2;
output 	MonDReg_23;
input 	writedata_23;
input 	writedata_24;
input 	byteenable_3;
output 	MonDReg_25;
input 	writedata_25;
output 	MonDReg_26;
input 	writedata_26;
output 	MonDReg_11;
input 	writedata_11;
input 	byteenable_1;
output 	MonDReg_13;
input 	writedata_13;
input 	writedata_16;
input 	writedata_12;
input 	jdo_23;
input 	writedata_5;
input 	writedata_4;
output 	MonDReg_14;
input 	writedata_14;
output 	MonDReg_15;
input 	writedata_15;
input 	writedata_18;
output 	MonDReg_17;
input 	writedata_17;
output 	MonDReg_10;
input 	writedata_10;
output 	MonDReg_9;
input 	writedata_9;
input 	writedata_8;
output 	MonDReg_7;
input 	writedata_7;
output 	MonDReg_6;
input 	writedata_6;
output 	MonDReg_21;
input 	writedata_21;
input 	writedata_19;
input 	writedata_20;
input 	jdo_16;
output 	MonDReg_31;
output 	MonDReg_30;
output 	MonDReg_28;
output 	MonDReg_27;
input 	jdo_7;
input 	jdo_24;
input 	jdo_22;
input 	jdo_14;
input 	jdo_15;
input 	jdo_8;
input 	writedata_27;
input 	writedata_28;
input 	writedata_29;
input 	writedata_30;
input 	writedata_31;
input 	jdo_13;
input 	jdo_12;
input 	jdo_11;
input 	jdo_10;
input 	jdo_9;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ociram_wr_en~0_combout ;
wire \jtag_ram_wr~q ;
wire \ociram_wr_en~1_combout ;
wire \ociram_reset_req~combout ;
wire \ociram_wr_data[0]~0_combout ;
wire \ociram_addr[0]~0_combout ;
wire \ociram_addr[1]~1_combout ;
wire \ociram_addr[2]~2_combout ;
wire \ociram_addr[3]~3_combout ;
wire \ociram_addr[4]~4_combout ;
wire \ociram_addr[5]~5_combout ;
wire \ociram_addr[6]~6_combout ;
wire \ociram_addr[7]~7_combout ;
wire \ociram_byteenable[0]~0_combout ;
wire \ociram_wr_data[1]~1_combout ;
wire \jtag_ram_wr~0_combout ;
wire \ociram_wr_data[2]~2_combout ;
wire \ociram_wr_data[22]~3_combout ;
wire \ociram_byteenable[2]~1_combout ;
wire \ociram_wr_data[23]~4_combout ;
wire \ociram_wr_data[24]~5_combout ;
wire \ociram_byteenable[3]~2_combout ;
wire \ociram_wr_data[25]~6_combout ;
wire \ociram_wr_data[26]~7_combout ;
wire \ociram_wr_data[11]~8_combout ;
wire \ociram_byteenable[1]~3_combout ;
wire \ociram_wr_data[13]~9_combout ;
wire \ociram_wr_data[16]~10_combout ;
wire \ociram_wr_data[12]~11_combout ;
wire \ociram_wr_data[3]~12_combout ;
wire \ociram_wr_data[5]~13_combout ;
wire \ociram_wr_data[4]~14_combout ;
wire \ociram_wr_data[14]~15_combout ;
wire \ociram_wr_data[15]~16_combout ;
wire \ociram_wr_data[18]~17_combout ;
wire \ociram_wr_data[17]~18_combout ;
wire \ociram_wr_data[10]~19_combout ;
wire \ociram_wr_data[9]~20_combout ;
wire \ociram_wr_data[8]~21_combout ;
wire \ociram_wr_data[7]~22_combout ;
wire \ociram_wr_data[6]~23_combout ;
wire \ociram_wr_data[21]~24_combout ;
wire \ociram_wr_data[19]~25_combout ;
wire \ociram_wr_data[20]~26_combout ;
wire \ociram_wr_data[27]~27_combout ;
wire \ociram_wr_data[28]~28_combout ;
wire \ociram_wr_data[29]~29_combout ;
wire \ociram_wr_data[30]~30_combout ;
wire \ociram_wr_data[31]~31_combout ;
wire \MonARegAddrInc[0]~0_combout ;
wire \MonAReg~7_combout ;
wire \MonAReg[2]~q ;
wire \MonARegAddrInc[0]~1 ;
wire \MonARegAddrInc[1]~2_combout ;
wire \MonAReg~6_combout ;
wire \MonAReg[3]~q ;
wire \MonARegAddrInc[1]~3 ;
wire \MonARegAddrInc[2]~4_combout ;
wire \MonAReg~5_combout ;
wire \MonAReg[4]~q ;
wire \Equal0~0_combout ;
wire \jtag_ram_access~0_combout ;
wire \MonAReg[10]~q ;
wire \MonARegAddrInc[2]~5 ;
wire \MonARegAddrInc[3]~6_combout ;
wire \MonAReg~4_combout ;
wire \MonAReg[5]~q ;
wire \MonARegAddrInc[3]~7 ;
wire \MonARegAddrInc[4]~8_combout ;
wire \MonAReg~3_combout ;
wire \MonAReg[6]~q ;
wire \MonARegAddrInc[4]~9 ;
wire \MonARegAddrInc[5]~10_combout ;
wire \MonAReg~2_combout ;
wire \MonAReg[7]~q ;
wire \MonARegAddrInc[5]~11 ;
wire \MonARegAddrInc[6]~12_combout ;
wire \MonAReg~1_combout ;
wire \MonAReg[8]~q ;
wire \MonARegAddrInc[6]~13 ;
wire \MonARegAddrInc[7]~14_combout ;
wire \MonAReg~0_combout ;
wire \MonAReg[9]~q ;
wire \MonARegAddrInc[7]~15 ;
wire \MonARegAddrInc[8]~16_combout ;
wire \jtag_ram_rd~0_combout ;
wire \jtag_ram_rd~1_combout ;
wire \jtag_ram_rd~q ;
wire \jtag_ram_rd_d1~q ;
wire \MonDReg[4]~0_combout ;
wire \jtag_rd~0_combout ;
wire \jtag_rd~q ;
wire \jtag_rd_d1~q ;
wire \MonDReg[0]~7_combout ;
wire \MonDReg[12]~2_combout ;
wire \Equal0~1_combout ;
wire \MonDReg[5]~1_combout ;
wire \Equal0~2_combout ;
wire \MonDReg[18]~3_combout ;
wire \Equal0~3_combout ;
wire \MonDReg[8]~4_combout ;
wire \Equal0~4_combout ;
wire \MonDReg[29]~5_combout ;
wire \jtag_ram_access~1_combout ;
wire \jtag_ram_access~q ;
wire \waitrequest~0_combout ;
wire \avalon_ociram_readdata_ready~0_combout ;
wire \avalon_ociram_readdata_ready~1_combout ;
wire \avalon_ociram_readdata_ready~q ;
wire \waitrequest~1_combout ;
wire \MonDReg~6_combout ;
wire \MonDReg~8_combout ;
wire \MonDReg~9_combout ;
wire \MonDReg~10_combout ;
wire \MonDReg~11_combout ;
wire \MonDReg~12_combout ;
wire \MonDReg~13_combout ;
wire \MonDReg~14_combout ;
wire \MonDReg~15_combout ;
wire \MonDReg~16_combout ;
wire \MonDReg~17_combout ;
wire \MonDReg~18_combout ;
wire \MonDReg~19_combout ;
wire \MonDReg~20_combout ;
wire \MonDReg~21_combout ;
wire \MonDReg~22_combout ;
wire \MonDReg~23_combout ;
wire \MonDReg~24_combout ;
wire \MonDReg~25_combout ;
wire \MonDReg~26_combout ;
wire \MonDReg~27_combout ;
wire \MonDReg~28_combout ;
wire \MonDReg~29_combout ;
wire \MonDReg~30_combout ;
wire \MonDReg~31_combout ;
wire \MonDReg~32_combout ;


nios_mcu_nios_mcu_nios_cpu_cpu_ociram_sp_ram_module nios_mcu_nios_cpu_cpu_ociram_sp_ram(
	.q_a_0(q_a_0),
	.q_a_1(q_a_1),
	.q_a_2(q_a_2),
	.q_a_22(q_a_22),
	.q_a_23(q_a_23),
	.q_a_24(q_a_24),
	.q_a_25(q_a_25),
	.q_a_26(q_a_26),
	.q_a_11(q_a_11),
	.q_a_13(q_a_13),
	.q_a_16(q_a_16),
	.q_a_12(q_a_12),
	.q_a_3(q_a_3),
	.q_a_5(q_a_5),
	.q_a_4(q_a_4),
	.q_a_14(q_a_14),
	.q_a_15(q_a_15),
	.q_a_18(q_a_18),
	.q_a_17(q_a_17),
	.q_a_10(q_a_10),
	.q_a_9(q_a_9),
	.q_a_8(q_a_8),
	.q_a_7(q_a_7),
	.q_a_6(q_a_6),
	.q_a_21(q_a_21),
	.q_a_19(q_a_19),
	.q_a_20(q_a_20),
	.q_a_27(q_a_27),
	.q_a_28(q_a_28),
	.q_a_29(q_a_29),
	.q_a_30(q_a_30),
	.q_a_31(q_a_31),
	.ociram_wr_en(\ociram_wr_en~1_combout ),
	.ociram_reset_req(\ociram_reset_req~combout ),
	.ociram_wr_data_0(\ociram_wr_data[0]~0_combout ),
	.ociram_addr_0(\ociram_addr[0]~0_combout ),
	.ociram_addr_1(\ociram_addr[1]~1_combout ),
	.ociram_addr_2(\ociram_addr[2]~2_combout ),
	.ociram_addr_3(\ociram_addr[3]~3_combout ),
	.ociram_addr_4(\ociram_addr[4]~4_combout ),
	.ociram_addr_5(\ociram_addr[5]~5_combout ),
	.ociram_addr_6(\ociram_addr[6]~6_combout ),
	.ociram_addr_7(\ociram_addr[7]~7_combout ),
	.ociram_byteenable_0(\ociram_byteenable[0]~0_combout ),
	.ociram_wr_data_1(\ociram_wr_data[1]~1_combout ),
	.ociram_wr_data_2(\ociram_wr_data[2]~2_combout ),
	.ociram_wr_data_22(\ociram_wr_data[22]~3_combout ),
	.ociram_byteenable_2(\ociram_byteenable[2]~1_combout ),
	.ociram_wr_data_23(\ociram_wr_data[23]~4_combout ),
	.ociram_wr_data_24(\ociram_wr_data[24]~5_combout ),
	.ociram_byteenable_3(\ociram_byteenable[3]~2_combout ),
	.ociram_wr_data_25(\ociram_wr_data[25]~6_combout ),
	.ociram_wr_data_26(\ociram_wr_data[26]~7_combout ),
	.ociram_wr_data_11(\ociram_wr_data[11]~8_combout ),
	.ociram_byteenable_1(\ociram_byteenable[1]~3_combout ),
	.ociram_wr_data_13(\ociram_wr_data[13]~9_combout ),
	.ociram_wr_data_16(\ociram_wr_data[16]~10_combout ),
	.ociram_wr_data_12(\ociram_wr_data[12]~11_combout ),
	.ociram_wr_data_3(\ociram_wr_data[3]~12_combout ),
	.ociram_wr_data_5(\ociram_wr_data[5]~13_combout ),
	.ociram_wr_data_4(\ociram_wr_data[4]~14_combout ),
	.ociram_wr_data_14(\ociram_wr_data[14]~15_combout ),
	.ociram_wr_data_15(\ociram_wr_data[15]~16_combout ),
	.ociram_wr_data_18(\ociram_wr_data[18]~17_combout ),
	.ociram_wr_data_17(\ociram_wr_data[17]~18_combout ),
	.ociram_wr_data_10(\ociram_wr_data[10]~19_combout ),
	.ociram_wr_data_9(\ociram_wr_data[9]~20_combout ),
	.ociram_wr_data_8(\ociram_wr_data[8]~21_combout ),
	.ociram_wr_data_7(\ociram_wr_data[7]~22_combout ),
	.ociram_wr_data_6(\ociram_wr_data[6]~23_combout ),
	.ociram_wr_data_21(\ociram_wr_data[21]~24_combout ),
	.ociram_wr_data_19(\ociram_wr_data[19]~25_combout ),
	.ociram_wr_data_20(\ociram_wr_data[20]~26_combout ),
	.ociram_wr_data_27(\ociram_wr_data[27]~27_combout ),
	.ociram_wr_data_28(\ociram_wr_data[28]~28_combout ),
	.ociram_wr_data_29(\ociram_wr_data[29]~29_combout ),
	.ociram_wr_data_30(\ociram_wr_data[30]~30_combout ),
	.ociram_wr_data_31(\ociram_wr_data[31]~31_combout ),
	.clk_clk(clk_clk));

cycloneive_lcell_comb \ociram_wr_en~0 (
	.dataa(write),
	.datab(debugaccess),
	.datac(address_8),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_en~0_combout ),
	.cout());
defparam \ociram_wr_en~0 .lut_mask = 16'hEFFF;
defparam \ociram_wr_en~0 .sum_lutc_input = "datac";

dffeas jtag_ram_wr(
	.clk(clk_clk),
	.d(\jtag_ram_wr~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_ram_wr~q ),
	.prn(vcc));
defparam jtag_ram_wr.is_wysiwyg = "true";
defparam jtag_ram_wr.power_up = "low";

cycloneive_lcell_comb \ociram_wr_en~1 (
	.dataa(\ociram_wr_en~0_combout ),
	.datab(\jtag_ram_access~q ),
	.datac(\jtag_ram_wr~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ociram_wr_en~1_combout ),
	.cout());
defparam \ociram_wr_en~1 .lut_mask = 16'hFEFE;
defparam \ociram_wr_en~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb ociram_reset_req(
	.dataa(r_early_rst),
	.datab(gnd),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_reset_req~combout ),
	.cout());
defparam ociram_reset_req.lut_mask = 16'hFF55;
defparam ociram_reset_req.sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[0]~0 (
	.dataa(MonDReg_0),
	.datab(writedata_0),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[0]~0_combout ),
	.cout());
defparam \ociram_wr_data[0]~0 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_addr[0]~0 (
	.dataa(\MonAReg[2]~q ),
	.datab(address_0),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[0]~0_combout ),
	.cout());
defparam \ociram_addr[0]~0 .lut_mask = 16'hAACC;
defparam \ociram_addr[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_addr[1]~1 (
	.dataa(\MonAReg[3]~q ),
	.datab(address_1),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[1]~1_combout ),
	.cout());
defparam \ociram_addr[1]~1 .lut_mask = 16'hAACC;
defparam \ociram_addr[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_addr[2]~2 (
	.dataa(\MonAReg[4]~q ),
	.datab(address_2),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[2]~2_combout ),
	.cout());
defparam \ociram_addr[2]~2 .lut_mask = 16'hAACC;
defparam \ociram_addr[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_addr[3]~3 (
	.dataa(\MonAReg[5]~q ),
	.datab(address_3),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[3]~3_combout ),
	.cout());
defparam \ociram_addr[3]~3 .lut_mask = 16'hAACC;
defparam \ociram_addr[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_addr[4]~4 (
	.dataa(\MonAReg[6]~q ),
	.datab(address_4),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[4]~4_combout ),
	.cout());
defparam \ociram_addr[4]~4 .lut_mask = 16'hAACC;
defparam \ociram_addr[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_addr[5]~5 (
	.dataa(\MonAReg[7]~q ),
	.datab(address_5),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[5]~5_combout ),
	.cout());
defparam \ociram_addr[5]~5 .lut_mask = 16'hAACC;
defparam \ociram_addr[5]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_addr[6]~6 (
	.dataa(\MonAReg[8]~q ),
	.datab(address_6),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[6]~6_combout ),
	.cout());
defparam \ociram_addr[6]~6 .lut_mask = 16'hAACC;
defparam \ociram_addr[6]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_addr[7]~7 (
	.dataa(\MonAReg[9]~q ),
	.datab(address_7),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_addr[7]~7_combout ),
	.cout());
defparam \ociram_addr[7]~7 .lut_mask = 16'hAACC;
defparam \ociram_addr[7]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_byteenable[0]~0 (
	.dataa(\jtag_ram_access~q ),
	.datab(byteenable_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ociram_byteenable[0]~0_combout ),
	.cout());
defparam \ociram_byteenable[0]~0 .lut_mask = 16'hEEEE;
defparam \ociram_byteenable[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[1]~1 (
	.dataa(MonDReg_1),
	.datab(writedata_1),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[1]~1_combout ),
	.cout());
defparam \ociram_wr_data[1]~1 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \jtag_ram_wr~0 (
	.dataa(take_action_ocimem_a),
	.datab(\jtag_ram_wr~q ),
	.datac(jdo_35),
	.datad(\MonARegAddrInc[8]~16_combout ),
	.cin(gnd),
	.combout(\jtag_ram_wr~0_combout ),
	.cout());
defparam \jtag_ram_wr~0 .lut_mask = 16'hACFF;
defparam \jtag_ram_wr~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[2]~2 (
	.dataa(MonDReg_2),
	.datab(writedata_2),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[2]~2_combout ),
	.cout());
defparam \ociram_wr_data[2]~2 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[22]~3 (
	.dataa(MonDReg_22),
	.datab(writedata_22),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[22]~3_combout ),
	.cout());
defparam \ociram_wr_data[22]~3 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[22]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_byteenable[2]~1 (
	.dataa(\jtag_ram_access~q ),
	.datab(byteenable_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ociram_byteenable[2]~1_combout ),
	.cout());
defparam \ociram_byteenable[2]~1 .lut_mask = 16'hEEEE;
defparam \ociram_byteenable[2]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[23]~4 (
	.dataa(MonDReg_23),
	.datab(writedata_23),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[23]~4_combout ),
	.cout());
defparam \ociram_wr_data[23]~4 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[23]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[24]~5 (
	.dataa(MonDReg_24),
	.datab(writedata_24),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[24]~5_combout ),
	.cout());
defparam \ociram_wr_data[24]~5 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[24]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_byteenable[3]~2 (
	.dataa(\jtag_ram_access~q ),
	.datab(byteenable_3),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ociram_byteenable[3]~2_combout ),
	.cout());
defparam \ociram_byteenable[3]~2 .lut_mask = 16'hEEEE;
defparam \ociram_byteenable[3]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[25]~6 (
	.dataa(MonDReg_25),
	.datab(writedata_25),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[25]~6_combout ),
	.cout());
defparam \ociram_wr_data[25]~6 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[25]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[26]~7 (
	.dataa(MonDReg_26),
	.datab(writedata_26),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[26]~7_combout ),
	.cout());
defparam \ociram_wr_data[26]~7 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[26]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[11]~8 (
	.dataa(MonDReg_11),
	.datab(writedata_11),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[11]~8_combout ),
	.cout());
defparam \ociram_wr_data[11]~8 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[11]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_byteenable[1]~3 (
	.dataa(\jtag_ram_access~q ),
	.datab(byteenable_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ociram_byteenable[1]~3_combout ),
	.cout());
defparam \ociram_byteenable[1]~3 .lut_mask = 16'hEEEE;
defparam \ociram_byteenable[1]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[13]~9 (
	.dataa(MonDReg_13),
	.datab(writedata_13),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[13]~9_combout ),
	.cout());
defparam \ociram_wr_data[13]~9 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[13]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[16]~10 (
	.dataa(MonDReg_16),
	.datab(writedata_16),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[16]~10_combout ),
	.cout());
defparam \ociram_wr_data[16]~10 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[16]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[12]~11 (
	.dataa(MonDReg_12),
	.datab(writedata_12),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[12]~11_combout ),
	.cout());
defparam \ociram_wr_data[12]~11 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[12]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[3]~12 (
	.dataa(MonDReg_3),
	.datab(writedata_3),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[3]~12_combout ),
	.cout());
defparam \ociram_wr_data[3]~12 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[3]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[5]~13 (
	.dataa(MonDReg_5),
	.datab(writedata_5),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[5]~13_combout ),
	.cout());
defparam \ociram_wr_data[5]~13 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[5]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[4]~14 (
	.dataa(MonDReg_4),
	.datab(writedata_4),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[4]~14_combout ),
	.cout());
defparam \ociram_wr_data[4]~14 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[4]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[14]~15 (
	.dataa(MonDReg_14),
	.datab(writedata_14),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[14]~15_combout ),
	.cout());
defparam \ociram_wr_data[14]~15 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[14]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[15]~16 (
	.dataa(MonDReg_15),
	.datab(writedata_15),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[15]~16_combout ),
	.cout());
defparam \ociram_wr_data[15]~16 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[15]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[18]~17 (
	.dataa(MonDReg_18),
	.datab(writedata_18),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[18]~17_combout ),
	.cout());
defparam \ociram_wr_data[18]~17 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[18]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[17]~18 (
	.dataa(MonDReg_17),
	.datab(writedata_17),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[17]~18_combout ),
	.cout());
defparam \ociram_wr_data[17]~18 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[17]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[10]~19 (
	.dataa(MonDReg_10),
	.datab(writedata_10),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[10]~19_combout ),
	.cout());
defparam \ociram_wr_data[10]~19 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[10]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[9]~20 (
	.dataa(MonDReg_9),
	.datab(writedata_9),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[9]~20_combout ),
	.cout());
defparam \ociram_wr_data[9]~20 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[9]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[8]~21 (
	.dataa(MonDReg_8),
	.datab(writedata_8),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[8]~21_combout ),
	.cout());
defparam \ociram_wr_data[8]~21 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[8]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[7]~22 (
	.dataa(MonDReg_7),
	.datab(writedata_7),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[7]~22_combout ),
	.cout());
defparam \ociram_wr_data[7]~22 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[7]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[6]~23 (
	.dataa(MonDReg_6),
	.datab(writedata_6),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[6]~23_combout ),
	.cout());
defparam \ociram_wr_data[6]~23 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[6]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[21]~24 (
	.dataa(MonDReg_21),
	.datab(writedata_21),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[21]~24_combout ),
	.cout());
defparam \ociram_wr_data[21]~24 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[21]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[19]~25 (
	.dataa(MonDReg_19),
	.datab(writedata_19),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[19]~25_combout ),
	.cout());
defparam \ociram_wr_data[19]~25 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[19]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[20]~26 (
	.dataa(MonDReg_20),
	.datab(writedata_20),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[20]~26_combout ),
	.cout());
defparam \ociram_wr_data[20]~26 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[20]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[27]~27 (
	.dataa(MonDReg_27),
	.datab(writedata_27),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[27]~27_combout ),
	.cout());
defparam \ociram_wr_data[27]~27 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[27]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[28]~28 (
	.dataa(MonDReg_28),
	.datab(writedata_28),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[28]~28_combout ),
	.cout());
defparam \ociram_wr_data[28]~28 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[28]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[29]~29 (
	.dataa(MonDReg_29),
	.datab(writedata_29),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[29]~29_combout ),
	.cout());
defparam \ociram_wr_data[29]~29 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[29]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[30]~30 (
	.dataa(MonDReg_30),
	.datab(writedata_30),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[30]~30_combout ),
	.cout());
defparam \ociram_wr_data[30]~30 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[30]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ociram_wr_data[31]~31 (
	.dataa(MonDReg_31),
	.datab(writedata_31),
	.datac(gnd),
	.datad(\jtag_ram_access~q ),
	.cin(gnd),
	.combout(\ociram_wr_data[31]~31_combout ),
	.cout());
defparam \ociram_wr_data[31]~31 .lut_mask = 16'hAACC;
defparam \ociram_wr_data[31]~31 .sum_lutc_input = "datac";

dffeas \MonDReg[4] (
	.clk(clk_clk),
	.d(\MonDReg[4]~0_combout ),
	.asdata(jdo_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~7_combout ),
	.q(MonDReg_4),
	.prn(vcc));
defparam \MonDReg[4] .is_wysiwyg = "true";
defparam \MonDReg[4] .power_up = "low";

dffeas \MonDReg[12] (
	.clk(clk_clk),
	.d(\MonDReg[12]~2_combout ),
	.asdata(jdo_15),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~7_combout ),
	.q(MonDReg_12),
	.prn(vcc));
defparam \MonDReg[12] .is_wysiwyg = "true";
defparam \MonDReg[12] .power_up = "low";

dffeas \MonDReg[5] (
	.clk(clk_clk),
	.d(\MonDReg[5]~1_combout ),
	.asdata(jdo_8),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~7_combout ),
	.q(MonDReg_5),
	.prn(vcc));
defparam \MonDReg[5] .is_wysiwyg = "true";
defparam \MonDReg[5] .power_up = "low";

dffeas \MonDReg[18] (
	.clk(clk_clk),
	.d(\MonDReg[18]~3_combout ),
	.asdata(jdo_21),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~7_combout ),
	.q(MonDReg_18),
	.prn(vcc));
defparam \MonDReg[18] .is_wysiwyg = "true";
defparam \MonDReg[18] .power_up = "low";

dffeas \MonDReg[8] (
	.clk(clk_clk),
	.d(\MonDReg[8]~4_combout ),
	.asdata(jdo_11),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~7_combout ),
	.q(MonDReg_8),
	.prn(vcc));
defparam \MonDReg[8] .is_wysiwyg = "true";
defparam \MonDReg[8] .power_up = "low";

dffeas \MonDReg[29] (
	.clk(clk_clk),
	.d(\MonDReg[29]~5_combout ),
	.asdata(jdo_32),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_b),
	.ena(\MonDReg[0]~7_combout ),
	.q(MonDReg_29),
	.prn(vcc));
defparam \MonDReg[29] .is_wysiwyg = "true";
defparam \MonDReg[29] .power_up = "low";

dffeas waitrequest(
	.clk(clk_clk),
	.d(\waitrequest~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(waitrequest1),
	.prn(vcc));
defparam waitrequest.is_wysiwyg = "true";
defparam waitrequest.power_up = "low";

dffeas \MonDReg[0] (
	.clk(clk_clk),
	.d(\MonDReg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~7_combout ),
	.q(MonDReg_0),
	.prn(vcc));
defparam \MonDReg[0] .is_wysiwyg = "true";
defparam \MonDReg[0] .power_up = "low";

dffeas \MonDReg[1] (
	.clk(clk_clk),
	.d(\MonDReg~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~7_combout ),
	.q(MonDReg_1),
	.prn(vcc));
defparam \MonDReg[1] .is_wysiwyg = "true";
defparam \MonDReg[1] .power_up = "low";

dffeas \MonDReg[2] (
	.clk(clk_clk),
	.d(\MonDReg~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~7_combout ),
	.q(MonDReg_2),
	.prn(vcc));
defparam \MonDReg[2] .is_wysiwyg = "true";
defparam \MonDReg[2] .power_up = "low";

dffeas \MonDReg[3] (
	.clk(clk_clk),
	.d(\MonDReg~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~7_combout ),
	.q(MonDReg_3),
	.prn(vcc));
defparam \MonDReg[3] .is_wysiwyg = "true";
defparam \MonDReg[3] .power_up = "low";

dffeas \MonDReg[16] (
	.clk(clk_clk),
	.d(\MonDReg~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~7_combout ),
	.q(MonDReg_16),
	.prn(vcc));
defparam \MonDReg[16] .is_wysiwyg = "true";
defparam \MonDReg[16] .power_up = "low";

dffeas \MonDReg[24] (
	.clk(clk_clk),
	.d(\MonDReg~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~7_combout ),
	.q(MonDReg_24),
	.prn(vcc));
defparam \MonDReg[24] .is_wysiwyg = "true";
defparam \MonDReg[24] .power_up = "low";

dffeas \MonDReg[20] (
	.clk(clk_clk),
	.d(\MonDReg~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~7_combout ),
	.q(MonDReg_20),
	.prn(vcc));
defparam \MonDReg[20] .is_wysiwyg = "true";
defparam \MonDReg[20] .power_up = "low";

dffeas \MonDReg[19] (
	.clk(clk_clk),
	.d(\MonDReg~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~7_combout ),
	.q(MonDReg_19),
	.prn(vcc));
defparam \MonDReg[19] .is_wysiwyg = "true";
defparam \MonDReg[19] .power_up = "low";

dffeas \MonDReg[22] (
	.clk(clk_clk),
	.d(\MonDReg~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~7_combout ),
	.q(MonDReg_22),
	.prn(vcc));
defparam \MonDReg[22] .is_wysiwyg = "true";
defparam \MonDReg[22] .power_up = "low";

dffeas \MonDReg[23] (
	.clk(clk_clk),
	.d(\MonDReg~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~7_combout ),
	.q(MonDReg_23),
	.prn(vcc));
defparam \MonDReg[23] .is_wysiwyg = "true";
defparam \MonDReg[23] .power_up = "low";

dffeas \MonDReg[25] (
	.clk(clk_clk),
	.d(\MonDReg~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~7_combout ),
	.q(MonDReg_25),
	.prn(vcc));
defparam \MonDReg[25] .is_wysiwyg = "true";
defparam \MonDReg[25] .power_up = "low";

dffeas \MonDReg[26] (
	.clk(clk_clk),
	.d(\MonDReg~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~7_combout ),
	.q(MonDReg_26),
	.prn(vcc));
defparam \MonDReg[26] .is_wysiwyg = "true";
defparam \MonDReg[26] .power_up = "low";

dffeas \MonDReg[11] (
	.clk(clk_clk),
	.d(\MonDReg~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~7_combout ),
	.q(MonDReg_11),
	.prn(vcc));
defparam \MonDReg[11] .is_wysiwyg = "true";
defparam \MonDReg[11] .power_up = "low";

dffeas \MonDReg[13] (
	.clk(clk_clk),
	.d(\MonDReg~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~7_combout ),
	.q(MonDReg_13),
	.prn(vcc));
defparam \MonDReg[13] .is_wysiwyg = "true";
defparam \MonDReg[13] .power_up = "low";

dffeas \MonDReg[14] (
	.clk(clk_clk),
	.d(\MonDReg~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~7_combout ),
	.q(MonDReg_14),
	.prn(vcc));
defparam \MonDReg[14] .is_wysiwyg = "true";
defparam \MonDReg[14] .power_up = "low";

dffeas \MonDReg[15] (
	.clk(clk_clk),
	.d(\MonDReg~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~7_combout ),
	.q(MonDReg_15),
	.prn(vcc));
defparam \MonDReg[15] .is_wysiwyg = "true";
defparam \MonDReg[15] .power_up = "low";

dffeas \MonDReg[17] (
	.clk(clk_clk),
	.d(\MonDReg~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~7_combout ),
	.q(MonDReg_17),
	.prn(vcc));
defparam \MonDReg[17] .is_wysiwyg = "true";
defparam \MonDReg[17] .power_up = "low";

dffeas \MonDReg[10] (
	.clk(clk_clk),
	.d(\MonDReg~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~7_combout ),
	.q(MonDReg_10),
	.prn(vcc));
defparam \MonDReg[10] .is_wysiwyg = "true";
defparam \MonDReg[10] .power_up = "low";

dffeas \MonDReg[9] (
	.clk(clk_clk),
	.d(\MonDReg~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~7_combout ),
	.q(MonDReg_9),
	.prn(vcc));
defparam \MonDReg[9] .is_wysiwyg = "true";
defparam \MonDReg[9] .power_up = "low";

dffeas \MonDReg[7] (
	.clk(clk_clk),
	.d(\MonDReg~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~7_combout ),
	.q(MonDReg_7),
	.prn(vcc));
defparam \MonDReg[7] .is_wysiwyg = "true";
defparam \MonDReg[7] .power_up = "low";

dffeas \MonDReg[6] (
	.clk(clk_clk),
	.d(\MonDReg~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~7_combout ),
	.q(MonDReg_6),
	.prn(vcc));
defparam \MonDReg[6] .is_wysiwyg = "true";
defparam \MonDReg[6] .power_up = "low";

dffeas \MonDReg[21] (
	.clk(clk_clk),
	.d(\MonDReg~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~7_combout ),
	.q(MonDReg_21),
	.prn(vcc));
defparam \MonDReg[21] .is_wysiwyg = "true";
defparam \MonDReg[21] .power_up = "low";

dffeas \MonDReg[31] (
	.clk(clk_clk),
	.d(\MonDReg~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~7_combout ),
	.q(MonDReg_31),
	.prn(vcc));
defparam \MonDReg[31] .is_wysiwyg = "true";
defparam \MonDReg[31] .power_up = "low";

dffeas \MonDReg[30] (
	.clk(clk_clk),
	.d(\MonDReg~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~7_combout ),
	.q(MonDReg_30),
	.prn(vcc));
defparam \MonDReg[30] .is_wysiwyg = "true";
defparam \MonDReg[30] .power_up = "low";

dffeas \MonDReg[28] (
	.clk(clk_clk),
	.d(\MonDReg~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~7_combout ),
	.q(MonDReg_28),
	.prn(vcc));
defparam \MonDReg[28] .is_wysiwyg = "true";
defparam \MonDReg[28] .power_up = "low";

dffeas \MonDReg[27] (
	.clk(clk_clk),
	.d(\MonDReg~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~7_combout ),
	.q(MonDReg_27),
	.prn(vcc));
defparam \MonDReg[27] .is_wysiwyg = "true";
defparam \MonDReg[27] .power_up = "low";

cycloneive_lcell_comb \MonARegAddrInc[0]~0 (
	.dataa(\MonAReg[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\MonARegAddrInc[0]~0_combout ),
	.cout(\MonARegAddrInc[0]~1 ));
defparam \MonARegAddrInc[0]~0 .lut_mask = 16'h55AA;
defparam \MonARegAddrInc[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonAReg~7 (
	.dataa(jdo_26),
	.datab(\MonARegAddrInc[0]~0_combout ),
	.datac(take_action_ocimem_a1),
	.datad(jdo_34),
	.cin(gnd),
	.combout(\MonAReg~7_combout ),
	.cout());
defparam \MonAReg~7 .lut_mask = 16'hEFFE;
defparam \MonAReg~7 .sum_lutc_input = "datac";

dffeas \MonAReg[2] (
	.clk(clk_clk),
	.d(\MonAReg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[2]~q ),
	.prn(vcc));
defparam \MonAReg[2] .is_wysiwyg = "true";
defparam \MonAReg[2] .power_up = "low";

cycloneive_lcell_comb \MonARegAddrInc[1]~2 (
	.dataa(\MonAReg[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\MonARegAddrInc[0]~1 ),
	.combout(\MonARegAddrInc[1]~2_combout ),
	.cout(\MonARegAddrInc[1]~3 ));
defparam \MonARegAddrInc[1]~2 .lut_mask = 16'h5A5F;
defparam \MonARegAddrInc[1]~2 .sum_lutc_input = "cin";

cycloneive_lcell_comb \MonAReg~6 (
	.dataa(jdo_27),
	.datab(\MonARegAddrInc[1]~2_combout ),
	.datac(take_action_ocimem_a1),
	.datad(jdo_34),
	.cin(gnd),
	.combout(\MonAReg~6_combout ),
	.cout());
defparam \MonAReg~6 .lut_mask = 16'hEFFE;
defparam \MonAReg~6 .sum_lutc_input = "datac";

dffeas \MonAReg[3] (
	.clk(clk_clk),
	.d(\MonAReg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[3]~q ),
	.prn(vcc));
defparam \MonAReg[3] .is_wysiwyg = "true";
defparam \MonAReg[3] .power_up = "low";

cycloneive_lcell_comb \MonARegAddrInc[2]~4 (
	.dataa(\MonAReg[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\MonARegAddrInc[1]~3 ),
	.combout(\MonARegAddrInc[2]~4_combout ),
	.cout(\MonARegAddrInc[2]~5 ));
defparam \MonARegAddrInc[2]~4 .lut_mask = 16'h5AAF;
defparam \MonARegAddrInc[2]~4 .sum_lutc_input = "cin";

cycloneive_lcell_comb \MonAReg~5 (
	.dataa(jdo_28),
	.datab(\MonARegAddrInc[2]~4_combout ),
	.datac(take_action_ocimem_a1),
	.datad(jdo_34),
	.cin(gnd),
	.combout(\MonAReg~5_combout ),
	.cout());
defparam \MonAReg~5 .lut_mask = 16'hEFFE;
defparam \MonAReg~5 .sum_lutc_input = "datac";

dffeas \MonAReg[4] (
	.clk(clk_clk),
	.d(\MonAReg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[4]~q ),
	.prn(vcc));
defparam \MonAReg[4] .is_wysiwyg = "true";
defparam \MonAReg[4] .power_up = "low";

cycloneive_lcell_comb \Equal0~0 (
	.dataa(\MonAReg[2]~q ),
	.datab(gnd),
	.datac(\MonAReg[4]~q ),
	.datad(\MonAReg[3]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hAFFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \jtag_ram_access~0 (
	.dataa(jdo_17),
	.datab(\MonARegAddrInc[8]~16_combout ),
	.datac(take_action_ocimem_a1),
	.datad(jdo_34),
	.cin(gnd),
	.combout(\jtag_ram_access~0_combout ),
	.cout());
defparam \jtag_ram_access~0 .lut_mask = 16'hEFFE;
defparam \jtag_ram_access~0 .sum_lutc_input = "datac";

dffeas \MonAReg[10] (
	.clk(clk_clk),
	.d(\jtag_ram_access~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[10]~q ),
	.prn(vcc));
defparam \MonAReg[10] .is_wysiwyg = "true";
defparam \MonAReg[10] .power_up = "low";

cycloneive_lcell_comb \MonARegAddrInc[3]~6 (
	.dataa(\MonAReg[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\MonARegAddrInc[2]~5 ),
	.combout(\MonARegAddrInc[3]~6_combout ),
	.cout(\MonARegAddrInc[3]~7 ));
defparam \MonARegAddrInc[3]~6 .lut_mask = 16'h5A5F;
defparam \MonARegAddrInc[3]~6 .sum_lutc_input = "cin";

cycloneive_lcell_comb \MonAReg~4 (
	.dataa(jdo_29),
	.datab(\MonARegAddrInc[3]~6_combout ),
	.datac(take_action_ocimem_a1),
	.datad(jdo_34),
	.cin(gnd),
	.combout(\MonAReg~4_combout ),
	.cout());
defparam \MonAReg~4 .lut_mask = 16'hEFFE;
defparam \MonAReg~4 .sum_lutc_input = "datac";

dffeas \MonAReg[5] (
	.clk(clk_clk),
	.d(\MonAReg~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[5]~q ),
	.prn(vcc));
defparam \MonAReg[5] .is_wysiwyg = "true";
defparam \MonAReg[5] .power_up = "low";

cycloneive_lcell_comb \MonARegAddrInc[4]~8 (
	.dataa(\MonAReg[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\MonARegAddrInc[3]~7 ),
	.combout(\MonARegAddrInc[4]~8_combout ),
	.cout(\MonARegAddrInc[4]~9 ));
defparam \MonARegAddrInc[4]~8 .lut_mask = 16'h5AAF;
defparam \MonARegAddrInc[4]~8 .sum_lutc_input = "cin";

cycloneive_lcell_comb \MonAReg~3 (
	.dataa(jdo_30),
	.datab(\MonARegAddrInc[4]~8_combout ),
	.datac(take_action_ocimem_a1),
	.datad(jdo_34),
	.cin(gnd),
	.combout(\MonAReg~3_combout ),
	.cout());
defparam \MonAReg~3 .lut_mask = 16'hEFFE;
defparam \MonAReg~3 .sum_lutc_input = "datac";

dffeas \MonAReg[6] (
	.clk(clk_clk),
	.d(\MonAReg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[6]~q ),
	.prn(vcc));
defparam \MonAReg[6] .is_wysiwyg = "true";
defparam \MonAReg[6] .power_up = "low";

cycloneive_lcell_comb \MonARegAddrInc[5]~10 (
	.dataa(\MonAReg[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\MonARegAddrInc[4]~9 ),
	.combout(\MonARegAddrInc[5]~10_combout ),
	.cout(\MonARegAddrInc[5]~11 ));
defparam \MonARegAddrInc[5]~10 .lut_mask = 16'h5A5F;
defparam \MonARegAddrInc[5]~10 .sum_lutc_input = "cin";

cycloneive_lcell_comb \MonAReg~2 (
	.dataa(jdo_31),
	.datab(\MonARegAddrInc[5]~10_combout ),
	.datac(take_action_ocimem_a1),
	.datad(jdo_34),
	.cin(gnd),
	.combout(\MonAReg~2_combout ),
	.cout());
defparam \MonAReg~2 .lut_mask = 16'hEFFE;
defparam \MonAReg~2 .sum_lutc_input = "datac";

dffeas \MonAReg[7] (
	.clk(clk_clk),
	.d(\MonAReg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[7]~q ),
	.prn(vcc));
defparam \MonAReg[7] .is_wysiwyg = "true";
defparam \MonAReg[7] .power_up = "low";

cycloneive_lcell_comb \MonARegAddrInc[6]~12 (
	.dataa(\MonAReg[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\MonARegAddrInc[5]~11 ),
	.combout(\MonARegAddrInc[6]~12_combout ),
	.cout(\MonARegAddrInc[6]~13 ));
defparam \MonARegAddrInc[6]~12 .lut_mask = 16'h5AAF;
defparam \MonARegAddrInc[6]~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \MonAReg~1 (
	.dataa(jdo_32),
	.datab(\MonARegAddrInc[6]~12_combout ),
	.datac(take_action_ocimem_a1),
	.datad(jdo_34),
	.cin(gnd),
	.combout(\MonAReg~1_combout ),
	.cout());
defparam \MonAReg~1 .lut_mask = 16'hEFFE;
defparam \MonAReg~1 .sum_lutc_input = "datac";

dffeas \MonAReg[8] (
	.clk(clk_clk),
	.d(\MonAReg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[8]~q ),
	.prn(vcc));
defparam \MonAReg[8] .is_wysiwyg = "true";
defparam \MonAReg[8] .power_up = "low";

cycloneive_lcell_comb \MonARegAddrInc[7]~14 (
	.dataa(\MonAReg[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\MonARegAddrInc[6]~13 ),
	.combout(\MonARegAddrInc[7]~14_combout ),
	.cout(\MonARegAddrInc[7]~15 ));
defparam \MonARegAddrInc[7]~14 .lut_mask = 16'h5A5F;
defparam \MonARegAddrInc[7]~14 .sum_lutc_input = "cin";

cycloneive_lcell_comb \MonAReg~0 (
	.dataa(jdo_33),
	.datab(\MonARegAddrInc[7]~14_combout ),
	.datac(take_action_ocimem_a1),
	.datad(jdo_34),
	.cin(gnd),
	.combout(\MonAReg~0_combout ),
	.cout());
defparam \MonAReg~0 .lut_mask = 16'hEFFE;
defparam \MonAReg~0 .sum_lutc_input = "datac";

dffeas \MonAReg[9] (
	.clk(clk_clk),
	.d(\MonAReg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[9]~q ),
	.prn(vcc));
defparam \MonAReg[9] .is_wysiwyg = "true";
defparam \MonAReg[9] .power_up = "low";

cycloneive_lcell_comb \MonARegAddrInc[8]~16 (
	.dataa(\MonAReg[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\MonARegAddrInc[7]~15 ),
	.combout(\MonARegAddrInc[8]~16_combout ),
	.cout());
defparam \MonARegAddrInc[8]~16 .lut_mask = 16'h5A5A;
defparam \MonARegAddrInc[8]~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \jtag_ram_rd~0 (
	.dataa(take_action_ocimem_a1),
	.datab(jdo_34),
	.datac(\MonARegAddrInc[8]~16_combout ),
	.datad(jdo_17),
	.cin(gnd),
	.combout(\jtag_ram_rd~0_combout ),
	.cout());
defparam \jtag_ram_rd~0 .lut_mask = 16'h8BFF;
defparam \jtag_ram_rd~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \jtag_ram_rd~1 (
	.dataa(\jtag_ram_rd~0_combout ),
	.datab(take_action_ocimem_b),
	.datac(\jtag_ram_rd~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\jtag_ram_rd~1_combout ),
	.cout());
defparam \jtag_ram_rd~1 .lut_mask = 16'hFEFE;
defparam \jtag_ram_rd~1 .sum_lutc_input = "datac";

dffeas jtag_ram_rd(
	.clk(clk_clk),
	.d(\jtag_ram_rd~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_ram_rd~q ),
	.prn(vcc));
defparam jtag_ram_rd.is_wysiwyg = "true";
defparam jtag_ram_rd.power_up = "low";

dffeas jtag_ram_rd_d1(
	.clk(clk_clk),
	.d(\jtag_ram_rd~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_ram_rd_d1~q ),
	.prn(vcc));
defparam jtag_ram_rd_d1.is_wysiwyg = "true";
defparam jtag_ram_rd_d1.power_up = "low";

cycloneive_lcell_comb \MonDReg[4]~0 (
	.dataa(\Equal0~0_combout ),
	.datab(q_a_4),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[4]~0_combout ),
	.cout());
defparam \MonDReg[4]~0 .lut_mask = 16'hAACC;
defparam \MonDReg[4]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \jtag_rd~0 (
	.dataa(take_action_ocimem_a),
	.datab(\jtag_rd~q ),
	.datac(gnd),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\jtag_rd~0_combout ),
	.cout());
defparam \jtag_rd~0 .lut_mask = 16'hEEFF;
defparam \jtag_rd~0 .sum_lutc_input = "datac";

dffeas jtag_rd(
	.clk(clk_clk),
	.d(\jtag_rd~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_rd~q ),
	.prn(vcc));
defparam jtag_rd.is_wysiwyg = "true";
defparam jtag_rd.power_up = "low";

dffeas jtag_rd_d1(
	.clk(clk_clk),
	.d(\jtag_rd~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_rd_d1~q ),
	.prn(vcc));
defparam jtag_rd_d1.is_wysiwyg = "true";
defparam jtag_rd_d1.power_up = "low";

cycloneive_lcell_comb \MonDReg[0]~7 (
	.dataa(gnd),
	.datab(take_action_ocimem_a),
	.datac(\jtag_rd_d1~q ),
	.datad(jdo_35),
	.cin(gnd),
	.combout(\MonDReg[0]~7_combout ),
	.cout());
defparam \MonDReg[0]~7 .lut_mask = 16'hF3C0;
defparam \MonDReg[0]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[12]~2 (
	.dataa(\Equal0~0_combout ),
	.datab(q_a_12),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[12]~2_combout ),
	.cout());
defparam \MonDReg[12]~2 .lut_mask = 16'hAACC;
defparam \MonDReg[12]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~1 (
	.dataa(gnd),
	.datab(\MonAReg[4]~q ),
	.datac(\MonAReg[3]~q ),
	.datad(\MonAReg[2]~q ),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'h3FFF;
defparam \Equal0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[5]~1 (
	.dataa(\Equal0~1_combout ),
	.datab(q_a_5),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[5]~1_combout ),
	.cout());
defparam \MonDReg[5]~1 .lut_mask = 16'hAACC;
defparam \MonDReg[5]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~2 (
	.dataa(\MonAReg[3]~q ),
	.datab(gnd),
	.datac(\MonAReg[4]~q ),
	.datad(\MonAReg[2]~q ),
	.cin(gnd),
	.combout(\Equal0~2_combout ),
	.cout());
defparam \Equal0~2 .lut_mask = 16'hAFFF;
defparam \Equal0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[18]~3 (
	.dataa(\Equal0~2_combout ),
	.datab(q_a_18),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[18]~3_combout ),
	.cout());
defparam \MonDReg[18]~3 .lut_mask = 16'hAACC;
defparam \MonDReg[18]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~3 (
	.dataa(\MonAReg[3]~q ),
	.datab(\MonAReg[2]~q ),
	.datac(gnd),
	.datad(\MonAReg[4]~q ),
	.cin(gnd),
	.combout(\Equal0~3_combout ),
	.cout());
defparam \Equal0~3 .lut_mask = 16'hEEFF;
defparam \Equal0~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[8]~4 (
	.dataa(\Equal0~3_combout ),
	.datab(q_a_8),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[8]~4_combout ),
	.cout());
defparam \MonDReg[8]~4 .lut_mask = 16'hAACC;
defparam \MonDReg[8]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~4 (
	.dataa(\MonAReg[4]~q ),
	.datab(gnd),
	.datac(\MonAReg[3]~q ),
	.datad(\MonAReg[2]~q ),
	.cin(gnd),
	.combout(\Equal0~4_combout ),
	.cout());
defparam \Equal0~4 .lut_mask = 16'hAFFF;
defparam \Equal0~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg[29]~5 (
	.dataa(\Equal0~4_combout ),
	.datab(q_a_29),
	.datac(gnd),
	.datad(\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.combout(\MonDReg[29]~5_combout ),
	.cout());
defparam \MonDReg[29]~5 .lut_mask = 16'hAACC;
defparam \MonDReg[29]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \jtag_ram_access~1 (
	.dataa(\jtag_ram_access~0_combout ),
	.datab(\MonARegAddrInc[8]~16_combout ),
	.datac(take_action_ocimem_b),
	.datad(take_action_ocimem_a1),
	.cin(gnd),
	.combout(\jtag_ram_access~1_combout ),
	.cout());
defparam \jtag_ram_access~1 .lut_mask = 16'hF377;
defparam \jtag_ram_access~1 .sum_lutc_input = "datac";

dffeas jtag_ram_access(
	.clk(clk_clk),
	.d(\jtag_ram_access~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_ram_access~q ),
	.prn(vcc));
defparam jtag_ram_access.is_wysiwyg = "true";
defparam jtag_ram_access.power_up = "low";

cycloneive_lcell_comb \waitrequest~0 (
	.dataa(write),
	.datab(\jtag_ram_access~q ),
	.datac(address_8),
	.datad(waitrequest1),
	.cin(gnd),
	.combout(\waitrequest~0_combout ),
	.cout());
defparam \waitrequest~0 .lut_mask = 16'hEFFF;
defparam \waitrequest~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \avalon_ociram_readdata_ready~0 (
	.dataa(read),
	.datab(address_8),
	.datac(\jtag_ram_access~q ),
	.datad(write),
	.cin(gnd),
	.combout(\avalon_ociram_readdata_ready~0_combout ),
	.cout());
defparam \avalon_ociram_readdata_ready~0 .lut_mask = 16'hEFFF;
defparam \avalon_ociram_readdata_ready~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \avalon_ociram_readdata_ready~1 (
	.dataa(waitrequest1),
	.datab(\avalon_ociram_readdata_ready~0_combout ),
	.datac(write),
	.datad(\avalon_ociram_readdata_ready~q ),
	.cin(gnd),
	.combout(\avalon_ociram_readdata_ready~1_combout ),
	.cout());
defparam \avalon_ociram_readdata_ready~1 .lut_mask = 16'hFFFE;
defparam \avalon_ociram_readdata_ready~1 .sum_lutc_input = "datac";

dffeas avalon_ociram_readdata_ready(
	.clk(clk_clk),
	.d(\avalon_ociram_readdata_ready~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\avalon_ociram_readdata_ready~q ),
	.prn(vcc));
defparam avalon_ociram_readdata_ready.is_wysiwyg = "true";
defparam avalon_ociram_readdata_ready.power_up = "low";

cycloneive_lcell_comb \waitrequest~1 (
	.dataa(\waitrequest~0_combout ),
	.datab(read),
	.datac(\avalon_ociram_readdata_ready~q ),
	.datad(write),
	.cin(gnd),
	.combout(\waitrequest~1_combout ),
	.cout());
defparam \waitrequest~1 .lut_mask = 16'hBFFF;
defparam \waitrequest~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~6 (
	.dataa(jdo_3),
	.datab(q_a_0),
	.datac(\jtag_ram_rd_d1~q ),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~6_combout ),
	.cout());
defparam \MonDReg~6 .lut_mask = 16'hFAFC;
defparam \MonDReg~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~8 (
	.dataa(jdo_4),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_1),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~8_combout ),
	.cout());
defparam \MonDReg~8 .lut_mask = 16'hFAFC;
defparam \MonDReg~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~9 (
	.dataa(jdo_5),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_2),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~9_combout ),
	.cout());
defparam \MonDReg~9 .lut_mask = 16'hFAFC;
defparam \MonDReg~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~10 (
	.dataa(jdo_6),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_3),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~10_combout ),
	.cout());
defparam \MonDReg~10 .lut_mask = 16'hFAFC;
defparam \MonDReg~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~11 (
	.dataa(jdo_19),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_16),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~11_combout ),
	.cout());
defparam \MonDReg~11 .lut_mask = 16'hFAFC;
defparam \MonDReg~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~12 (
	.dataa(jdo_27),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_24),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~12_combout ),
	.cout());
defparam \MonDReg~12 .lut_mask = 16'hFAFC;
defparam \MonDReg~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~13 (
	.dataa(jdo_23),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_20),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~13_combout ),
	.cout());
defparam \MonDReg~13 .lut_mask = 16'hFAFC;
defparam \MonDReg~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~14 (
	.dataa(jdo_22),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_19),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~14_combout ),
	.cout());
defparam \MonDReg~14 .lut_mask = 16'hFAFC;
defparam \MonDReg~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~15 (
	.dataa(jdo_25),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_22),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~15_combout ),
	.cout());
defparam \MonDReg~15 .lut_mask = 16'hFAFC;
defparam \MonDReg~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~16 (
	.dataa(jdo_26),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_23),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~16_combout ),
	.cout());
defparam \MonDReg~16 .lut_mask = 16'hFAFC;
defparam \MonDReg~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~17 (
	.dataa(jdo_28),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_25),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~17_combout ),
	.cout());
defparam \MonDReg~17 .lut_mask = 16'hFAFC;
defparam \MonDReg~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~18 (
	.dataa(jdo_29),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_26),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~18_combout ),
	.cout());
defparam \MonDReg~18 .lut_mask = 16'hFAFC;
defparam \MonDReg~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~19 (
	.dataa(jdo_14),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_11),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~19_combout ),
	.cout());
defparam \MonDReg~19 .lut_mask = 16'hFAFC;
defparam \MonDReg~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~20 (
	.dataa(jdo_16),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_13),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~20_combout ),
	.cout());
defparam \MonDReg~20 .lut_mask = 16'hFAFC;
defparam \MonDReg~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~21 (
	.dataa(jdo_17),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_14),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~21_combout ),
	.cout());
defparam \MonDReg~21 .lut_mask = 16'hFAFC;
defparam \MonDReg~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~22 (
	.dataa(jdo_18),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_15),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~22_combout ),
	.cout());
defparam \MonDReg~22 .lut_mask = 16'hFAFC;
defparam \MonDReg~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~23 (
	.dataa(jdo_20),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_17),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~23_combout ),
	.cout());
defparam \MonDReg~23 .lut_mask = 16'hFAFC;
defparam \MonDReg~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~24 (
	.dataa(jdo_13),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_10),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~24_combout ),
	.cout());
defparam \MonDReg~24 .lut_mask = 16'hFAFC;
defparam \MonDReg~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~25 (
	.dataa(jdo_12),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_9),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~25_combout ),
	.cout());
defparam \MonDReg~25 .lut_mask = 16'hFAFC;
defparam \MonDReg~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~26 (
	.dataa(jdo_10),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_7),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~26_combout ),
	.cout());
defparam \MonDReg~26 .lut_mask = 16'hFAFC;
defparam \MonDReg~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~27 (
	.dataa(jdo_9),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_6),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~27_combout ),
	.cout());
defparam \MonDReg~27 .lut_mask = 16'hFAFC;
defparam \MonDReg~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~28 (
	.dataa(jdo_24),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_21),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~28_combout ),
	.cout());
defparam \MonDReg~28 .lut_mask = 16'hFAFC;
defparam \MonDReg~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~29 (
	.dataa(jdo_34),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_31),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~29_combout ),
	.cout());
defparam \MonDReg~29 .lut_mask = 16'hFAFC;
defparam \MonDReg~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~30 (
	.dataa(jdo_33),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_30),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~30_combout ),
	.cout());
defparam \MonDReg~30 .lut_mask = 16'hFAFC;
defparam \MonDReg~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~31 (
	.dataa(jdo_31),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_28),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~31_combout ),
	.cout());
defparam \MonDReg~31 .lut_mask = 16'hFAFC;
defparam \MonDReg~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \MonDReg~32 (
	.dataa(jdo_30),
	.datab(\jtag_ram_rd_d1~q ),
	.datac(q_a_27),
	.datad(take_action_ocimem_b),
	.cin(gnd),
	.combout(\MonDReg~32_combout ),
	.cout());
defparam \MonDReg~32 .lut_mask = 16'hFAFC;
defparam \MonDReg~32 .sum_lutc_input = "datac";

endmodule

module nios_mcu_nios_mcu_nios_cpu_cpu_ociram_sp_ram_module (
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_22,
	q_a_23,
	q_a_24,
	q_a_25,
	q_a_26,
	q_a_11,
	q_a_13,
	q_a_16,
	q_a_12,
	q_a_3,
	q_a_5,
	q_a_4,
	q_a_14,
	q_a_15,
	q_a_18,
	q_a_17,
	q_a_10,
	q_a_9,
	q_a_8,
	q_a_7,
	q_a_6,
	q_a_21,
	q_a_19,
	q_a_20,
	q_a_27,
	q_a_28,
	q_a_29,
	q_a_30,
	q_a_31,
	ociram_wr_en,
	ociram_reset_req,
	ociram_wr_data_0,
	ociram_addr_0,
	ociram_addr_1,
	ociram_addr_2,
	ociram_addr_3,
	ociram_addr_4,
	ociram_addr_5,
	ociram_addr_6,
	ociram_addr_7,
	ociram_byteenable_0,
	ociram_wr_data_1,
	ociram_wr_data_2,
	ociram_wr_data_22,
	ociram_byteenable_2,
	ociram_wr_data_23,
	ociram_wr_data_24,
	ociram_byteenable_3,
	ociram_wr_data_25,
	ociram_wr_data_26,
	ociram_wr_data_11,
	ociram_byteenable_1,
	ociram_wr_data_13,
	ociram_wr_data_16,
	ociram_wr_data_12,
	ociram_wr_data_3,
	ociram_wr_data_5,
	ociram_wr_data_4,
	ociram_wr_data_14,
	ociram_wr_data_15,
	ociram_wr_data_18,
	ociram_wr_data_17,
	ociram_wr_data_10,
	ociram_wr_data_9,
	ociram_wr_data_8,
	ociram_wr_data_7,
	ociram_wr_data_6,
	ociram_wr_data_21,
	ociram_wr_data_19,
	ociram_wr_data_20,
	ociram_wr_data_27,
	ociram_wr_data_28,
	ociram_wr_data_29,
	ociram_wr_data_30,
	ociram_wr_data_31,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_22;
output 	q_a_23;
output 	q_a_24;
output 	q_a_25;
output 	q_a_26;
output 	q_a_11;
output 	q_a_13;
output 	q_a_16;
output 	q_a_12;
output 	q_a_3;
output 	q_a_5;
output 	q_a_4;
output 	q_a_14;
output 	q_a_15;
output 	q_a_18;
output 	q_a_17;
output 	q_a_10;
output 	q_a_9;
output 	q_a_8;
output 	q_a_7;
output 	q_a_6;
output 	q_a_21;
output 	q_a_19;
output 	q_a_20;
output 	q_a_27;
output 	q_a_28;
output 	q_a_29;
output 	q_a_30;
output 	q_a_31;
input 	ociram_wr_en;
input 	ociram_reset_req;
input 	ociram_wr_data_0;
input 	ociram_addr_0;
input 	ociram_addr_1;
input 	ociram_addr_2;
input 	ociram_addr_3;
input 	ociram_addr_4;
input 	ociram_addr_5;
input 	ociram_addr_6;
input 	ociram_addr_7;
input 	ociram_byteenable_0;
input 	ociram_wr_data_1;
input 	ociram_wr_data_2;
input 	ociram_wr_data_22;
input 	ociram_byteenable_2;
input 	ociram_wr_data_23;
input 	ociram_wr_data_24;
input 	ociram_byteenable_3;
input 	ociram_wr_data_25;
input 	ociram_wr_data_26;
input 	ociram_wr_data_11;
input 	ociram_byteenable_1;
input 	ociram_wr_data_13;
input 	ociram_wr_data_16;
input 	ociram_wr_data_12;
input 	ociram_wr_data_3;
input 	ociram_wr_data_5;
input 	ociram_wr_data_4;
input 	ociram_wr_data_14;
input 	ociram_wr_data_15;
input 	ociram_wr_data_18;
input 	ociram_wr_data_17;
input 	ociram_wr_data_10;
input 	ociram_wr_data_9;
input 	ociram_wr_data_8;
input 	ociram_wr_data_7;
input 	ociram_wr_data_6;
input 	ociram_wr_data_21;
input 	ociram_wr_data_19;
input 	ociram_wr_data_20;
input 	ociram_wr_data_27;
input 	ociram_wr_data_28;
input 	ociram_wr_data_29;
input 	ociram_wr_data_30;
input 	ociram_wr_data_31;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nios_mcu_altsyncram_1 the_altsyncram(
	.q_a({q_a_31,q_a_30,q_a_29,q_a_28,q_a_27,q_a_26,q_a_25,q_a_24,q_a_23,q_a_22,q_a_21,q_a_20,q_a_19,q_a_18,q_a_17,q_a_16,q_a_15,q_a_14,q_a_13,q_a_12,q_a_11,q_a_10,q_a_9,q_a_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.wren_a(ociram_wr_en),
	.clocken0(ociram_reset_req),
	.data_a({ociram_wr_data_31,ociram_wr_data_30,ociram_wr_data_29,ociram_wr_data_28,ociram_wr_data_27,ociram_wr_data_26,ociram_wr_data_25,ociram_wr_data_24,ociram_wr_data_23,ociram_wr_data_22,ociram_wr_data_21,ociram_wr_data_20,ociram_wr_data_19,ociram_wr_data_18,ociram_wr_data_17,
ociram_wr_data_16,ociram_wr_data_15,ociram_wr_data_14,ociram_wr_data_13,ociram_wr_data_12,ociram_wr_data_11,ociram_wr_data_10,ociram_wr_data_9,ociram_wr_data_8,ociram_wr_data_7,ociram_wr_data_6,ociram_wr_data_5,ociram_wr_data_4,ociram_wr_data_3,ociram_wr_data_2,
ociram_wr_data_1,ociram_wr_data_0}),
	.address_a({gnd,gnd,gnd,gnd,gnd,ociram_addr_7,ociram_addr_6,ociram_addr_5,ociram_addr_4,ociram_addr_3,ociram_addr_2,ociram_addr_1,ociram_addr_0}),
	.byteena_a({ociram_byteenable_3,ociram_byteenable_2,ociram_byteenable_1,ociram_byteenable_0}),
	.clock0(clk_clk));

endmodule

module nios_mcu_altsyncram_1 (
	q_a,
	wren_a,
	clocken0,
	data_a,
	address_a,
	byteena_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_a;
input 	wren_a;
input 	clocken0;
input 	[31:0] data_a;
input 	[12:0] address_a;
input 	[3:0] byteena_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nios_mcu_altsyncram_ac71 auto_generated(
	.q_a({q_a[31],q_a[30],q_a[29],q_a[28],q_a[27],q_a[26],q_a[25],q_a[24],q_a[23],q_a[22],q_a[21],q_a[20],q_a[19],q_a[18],q_a[17],q_a[16],q_a[15],q_a[14],q_a[13],q_a[12],q_a[11],q_a[10],q_a[9],q_a[8],q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.wren_a(wren_a),
	.clocken0(clocken0),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.byteena_a({byteena_a[3],byteena_a[2],byteena_a[1],byteena_a[0]}),
	.clock0(clock0));

endmodule

module nios_mcu_altsyncram_ac71 (
	q_a,
	wren_a,
	clocken0,
	data_a,
	address_a,
	byteena_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_a;
input 	wren_a;
input 	clocken0;
input 	[31:0] data_a;
input 	[7:0] address_a;
input 	[3:0] byteena_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a22_PORTADATAOUT_bus;
wire [143:0] ram_block1a23_PORTADATAOUT_bus;
wire [143:0] ram_block1a24_PORTADATAOUT_bus;
wire [143:0] ram_block1a25_PORTADATAOUT_bus;
wire [143:0] ram_block1a26_PORTADATAOUT_bus;
wire [143:0] ram_block1a11_PORTADATAOUT_bus;
wire [143:0] ram_block1a13_PORTADATAOUT_bus;
wire [143:0] ram_block1a16_PORTADATAOUT_bus;
wire [143:0] ram_block1a12_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a14_PORTADATAOUT_bus;
wire [143:0] ram_block1a15_PORTADATAOUT_bus;
wire [143:0] ram_block1a18_PORTADATAOUT_bus;
wire [143:0] ram_block1a17_PORTADATAOUT_bus;
wire [143:0] ram_block1a10_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a21_PORTADATAOUT_bus;
wire [143:0] ram_block1a19_PORTADATAOUT_bus;
wire [143:0] ram_block1a20_PORTADATAOUT_bus;
wire [143:0] ram_block1a27_PORTADATAOUT_bus;
wire [143:0] ram_block1a28_PORTADATAOUT_bus;
wire [143:0] ram_block1a29_PORTADATAOUT_bus;
wire [143:0] ram_block1a30_PORTADATAOUT_bus;
wire [143:0] ram_block1a31_PORTADATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[22] = ram_block1a22_PORTADATAOUT_bus[0];

assign q_a[23] = ram_block1a23_PORTADATAOUT_bus[0];

assign q_a[24] = ram_block1a24_PORTADATAOUT_bus[0];

assign q_a[25] = ram_block1a25_PORTADATAOUT_bus[0];

assign q_a[26] = ram_block1a26_PORTADATAOUT_bus[0];

assign q_a[11] = ram_block1a11_PORTADATAOUT_bus[0];

assign q_a[13] = ram_block1a13_PORTADATAOUT_bus[0];

assign q_a[16] = ram_block1a16_PORTADATAOUT_bus[0];

assign q_a[12] = ram_block1a12_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[14] = ram_block1a14_PORTADATAOUT_bus[0];

assign q_a[15] = ram_block1a15_PORTADATAOUT_bus[0];

assign q_a[18] = ram_block1a18_PORTADATAOUT_bus[0];

assign q_a[17] = ram_block1a17_PORTADATAOUT_bus[0];

assign q_a[10] = ram_block1a10_PORTADATAOUT_bus[0];

assign q_a[9] = ram_block1a9_PORTADATAOUT_bus[0];

assign q_a[8] = ram_block1a8_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[21] = ram_block1a21_PORTADATAOUT_bus[0];

assign q_a[19] = ram_block1a19_PORTADATAOUT_bus[0];

assign q_a[20] = ram_block1a20_PORTADATAOUT_bus[0];

assign q_a[27] = ram_block1a27_PORTADATAOUT_bus[0];

assign q_a[28] = ram_block1a28_PORTADATAOUT_bus[0];

assign q_a[29] = ram_block1a29_PORTADATAOUT_bus[0];

assign q_a[30] = ram_block1a30_PORTADATAOUT_bus[0];

assign q_a[31] = ram_block1a31_PORTADATAOUT_bus[0];

cycloneive_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_nios2_oci:the_nios_mcu_nios_cpu_cpu_nios2_oci|nios_mcu_nios_cpu_cpu_nios2_ocimem:the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram_module:nios_mcu_nios_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "single_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 8;
defparam ram_block1a0.port_a_byte_enable_mask_width = 1;
defparam ram_block1a0.port_a_byte_size = 1;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 255;
defparam ram_block1a0.port_a_logical_ram_depth = 256;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.ram_block_type = "auto";

cycloneive_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_nios2_oci:the_nios_mcu_nios_cpu_cpu_nios2_oci|nios_mcu_nios_cpu_cpu_nios2_ocimem:the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram_module:nios_mcu_nios_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "single_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 8;
defparam ram_block1a1.port_a_byte_enable_mask_width = 1;
defparam ram_block1a1.port_a_byte_size = 1;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 255;
defparam ram_block1a1.port_a_logical_ram_depth = 256;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.ram_block_type = "auto";

cycloneive_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_nios2_oci:the_nios_mcu_nios_cpu_cpu_nios2_oci|nios_mcu_nios_cpu_cpu_nios2_ocimem:the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram_module:nios_mcu_nios_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "single_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 8;
defparam ram_block1a2.port_a_byte_enable_mask_width = 1;
defparam ram_block1a2.port_a_byte_size = 1;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 255;
defparam ram_block1a2.port_a_logical_ram_depth = 256;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.ram_block_type = "auto";

cycloneive_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a22_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk0_input_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_nios2_oci:the_nios_mcu_nios_cpu_cpu_nios2_oci|nios_mcu_nios_cpu_cpu_nios2_ocimem:the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram_module:nios_mcu_nios_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.operation_mode = "single_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 8;
defparam ram_block1a22.port_a_byte_enable_mask_width = 1;
defparam ram_block1a22.port_a_byte_size = 1;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 255;
defparam ram_block1a22.port_a_logical_ram_depth = 256;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.ram_block_type = "auto";

cycloneive_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a23_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk0_input_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_nios2_oci:the_nios_mcu_nios_cpu_cpu_nios2_oci|nios_mcu_nios_cpu_cpu_nios2_ocimem:the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram_module:nios_mcu_nios_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.operation_mode = "single_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 8;
defparam ram_block1a23.port_a_byte_enable_mask_width = 1;
defparam ram_block1a23.port_a_byte_size = 1;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 255;
defparam ram_block1a23.port_a_logical_ram_depth = 256;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.ram_block_type = "auto";

cycloneive_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a24_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk0_input_clock_enable = "ena0";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_nios2_oci:the_nios_mcu_nios_cpu_cpu_nios2_oci|nios_mcu_nios_cpu_cpu_nios2_ocimem:the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram_module:nios_mcu_nios_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.operation_mode = "single_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 8;
defparam ram_block1a24.port_a_byte_enable_mask_width = 1;
defparam ram_block1a24.port_a_byte_size = 1;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 255;
defparam ram_block1a24.port_a_logical_ram_depth = 256;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.ram_block_type = "auto";

cycloneive_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a25_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk0_input_clock_enable = "ena0";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_nios2_oci:the_nios_mcu_nios_cpu_cpu_nios2_oci|nios_mcu_nios_cpu_cpu_nios2_ocimem:the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram_module:nios_mcu_nios_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.operation_mode = "single_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 8;
defparam ram_block1a25.port_a_byte_enable_mask_width = 1;
defparam ram_block1a25.port_a_byte_size = 1;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 255;
defparam ram_block1a25.port_a_logical_ram_depth = 256;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.ram_block_type = "auto";

cycloneive_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a26_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk0_input_clock_enable = "ena0";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_nios2_oci:the_nios_mcu_nios_cpu_cpu_nios2_oci|nios_mcu_nios_cpu_cpu_nios2_ocimem:the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram_module:nios_mcu_nios_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.operation_mode = "single_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 8;
defparam ram_block1a26.port_a_byte_enable_mask_width = 1;
defparam ram_block1a26.port_a_byte_size = 1;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 255;
defparam ram_block1a26.port_a_logical_ram_depth = 256;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a11_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_nios2_oci:the_nios_mcu_nios_cpu_cpu_nios2_oci|nios_mcu_nios_cpu_cpu_nios2_ocimem:the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram_module:nios_mcu_nios_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.operation_mode = "single_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 8;
defparam ram_block1a11.port_a_byte_enable_mask_width = 1;
defparam ram_block1a11.port_a_byte_size = 1;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 255;
defparam ram_block1a11.port_a_logical_ram_depth = 256;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a13_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_nios2_oci:the_nios_mcu_nios_cpu_cpu_nios2_oci|nios_mcu_nios_cpu_cpu_nios2_ocimem:the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram_module:nios_mcu_nios_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.operation_mode = "single_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 8;
defparam ram_block1a13.port_a_byte_enable_mask_width = 1;
defparam ram_block1a13.port_a_byte_size = 1;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 255;
defparam ram_block1a13.port_a_logical_ram_depth = 256;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a16_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_nios2_oci:the_nios_mcu_nios_cpu_cpu_nios2_oci|nios_mcu_nios_cpu_cpu_nios2_ocimem:the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram_module:nios_mcu_nios_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.operation_mode = "single_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 8;
defparam ram_block1a16.port_a_byte_enable_mask_width = 1;
defparam ram_block1a16.port_a_byte_size = 1;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 255;
defparam ram_block1a16.port_a_logical_ram_depth = 256;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a12_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_nios2_oci:the_nios_mcu_nios_cpu_cpu_nios2_oci|nios_mcu_nios_cpu_cpu_nios2_ocimem:the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram_module:nios_mcu_nios_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.operation_mode = "single_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 8;
defparam ram_block1a12.port_a_byte_enable_mask_width = 1;
defparam ram_block1a12.port_a_byte_size = 1;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 255;
defparam ram_block1a12.port_a_logical_ram_depth = 256;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_nios2_oci:the_nios_mcu_nios_cpu_cpu_nios2_oci|nios_mcu_nios_cpu_cpu_nios2_ocimem:the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram_module:nios_mcu_nios_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "single_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 8;
defparam ram_block1a3.port_a_byte_enable_mask_width = 1;
defparam ram_block1a3.port_a_byte_size = 1;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 255;
defparam ram_block1a3.port_a_logical_ram_depth = 256;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_nios2_oci:the_nios_mcu_nios_cpu_cpu_nios2_oci|nios_mcu_nios_cpu_cpu_nios2_ocimem:the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram_module:nios_mcu_nios_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "single_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 8;
defparam ram_block1a5.port_a_byte_enable_mask_width = 1;
defparam ram_block1a5.port_a_byte_size = 1;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 255;
defparam ram_block1a5.port_a_logical_ram_depth = 256;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_nios2_oci:the_nios_mcu_nios_cpu_cpu_nios2_oci|nios_mcu_nios_cpu_cpu_nios2_ocimem:the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram_module:nios_mcu_nios_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "single_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 8;
defparam ram_block1a4.port_a_byte_enable_mask_width = 1;
defparam ram_block1a4.port_a_byte_size = 1;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 255;
defparam ram_block1a4.port_a_logical_ram_depth = 256;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a14_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_nios2_oci:the_nios_mcu_nios_cpu_cpu_nios2_oci|nios_mcu_nios_cpu_cpu_nios2_ocimem:the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram_module:nios_mcu_nios_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.operation_mode = "single_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 8;
defparam ram_block1a14.port_a_byte_enable_mask_width = 1;
defparam ram_block1a14.port_a_byte_size = 1;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 255;
defparam ram_block1a14.port_a_logical_ram_depth = 256;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a15_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_nios2_oci:the_nios_mcu_nios_cpu_cpu_nios2_oci|nios_mcu_nios_cpu_cpu_nios2_ocimem:the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram_module:nios_mcu_nios_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.operation_mode = "single_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 8;
defparam ram_block1a15.port_a_byte_enable_mask_width = 1;
defparam ram_block1a15.port_a_byte_size = 1;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 255;
defparam ram_block1a15.port_a_logical_ram_depth = 256;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a18_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_nios2_oci:the_nios_mcu_nios_cpu_cpu_nios2_oci|nios_mcu_nios_cpu_cpu_nios2_ocimem:the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram_module:nios_mcu_nios_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.operation_mode = "single_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 8;
defparam ram_block1a18.port_a_byte_enable_mask_width = 1;
defparam ram_block1a18.port_a_byte_size = 1;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 255;
defparam ram_block1a18.port_a_logical_ram_depth = 256;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a17_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_nios2_oci:the_nios_mcu_nios_cpu_cpu_nios2_oci|nios_mcu_nios_cpu_cpu_nios2_ocimem:the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram_module:nios_mcu_nios_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.operation_mode = "single_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 8;
defparam ram_block1a17.port_a_byte_enable_mask_width = 1;
defparam ram_block1a17.port_a_byte_size = 1;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 255;
defparam ram_block1a17.port_a_logical_ram_depth = 256;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a10_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_nios2_oci:the_nios_mcu_nios_cpu_cpu_nios2_oci|nios_mcu_nios_cpu_cpu_nios2_ocimem:the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram_module:nios_mcu_nios_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.operation_mode = "single_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 8;
defparam ram_block1a10.port_a_byte_enable_mask_width = 1;
defparam ram_block1a10.port_a_byte_size = 1;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 255;
defparam ram_block1a10.port_a_logical_ram_depth = 256;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_nios2_oci:the_nios_mcu_nios_cpu_cpu_nios2_oci|nios_mcu_nios_cpu_cpu_nios2_ocimem:the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram_module:nios_mcu_nios_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.operation_mode = "single_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 8;
defparam ram_block1a9.port_a_byte_enable_mask_width = 1;
defparam ram_block1a9.port_a_byte_size = 1;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 255;
defparam ram_block1a9.port_a_logical_ram_depth = 256;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_nios2_oci:the_nios_mcu_nios_cpu_cpu_nios2_oci|nios_mcu_nios_cpu_cpu_nios2_ocimem:the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram_module:nios_mcu_nios_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.operation_mode = "single_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 8;
defparam ram_block1a8.port_a_byte_enable_mask_width = 1;
defparam ram_block1a8.port_a_byte_size = 1;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 255;
defparam ram_block1a8.port_a_logical_ram_depth = 256;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_nios2_oci:the_nios_mcu_nios_cpu_cpu_nios2_oci|nios_mcu_nios_cpu_cpu_nios2_ocimem:the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram_module:nios_mcu_nios_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "single_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 8;
defparam ram_block1a7.port_a_byte_enable_mask_width = 1;
defparam ram_block1a7.port_a_byte_size = 1;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 255;
defparam ram_block1a7.port_a_logical_ram_depth = 256;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_nios2_oci:the_nios_mcu_nios_cpu_cpu_nios2_oci|nios_mcu_nios_cpu_cpu_nios2_ocimem:the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram_module:nios_mcu_nios_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "single_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 8;
defparam ram_block1a6.port_a_byte_enable_mask_width = 1;
defparam ram_block1a6.port_a_byte_size = 1;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 255;
defparam ram_block1a6.port_a_logical_ram_depth = 256;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a21_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk0_input_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_nios2_oci:the_nios_mcu_nios_cpu_cpu_nios2_oci|nios_mcu_nios_cpu_cpu_nios2_ocimem:the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram_module:nios_mcu_nios_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.operation_mode = "single_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 8;
defparam ram_block1a21.port_a_byte_enable_mask_width = 1;
defparam ram_block1a21.port_a_byte_size = 1;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 255;
defparam ram_block1a21.port_a_logical_ram_depth = 256;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a19_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_nios2_oci:the_nios_mcu_nios_cpu_cpu_nios2_oci|nios_mcu_nios_cpu_cpu_nios2_ocimem:the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram_module:nios_mcu_nios_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.operation_mode = "single_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 8;
defparam ram_block1a19.port_a_byte_enable_mask_width = 1;
defparam ram_block1a19.port_a_byte_size = 1;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 255;
defparam ram_block1a19.port_a_logical_ram_depth = 256;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.ram_block_type = "auto";

cycloneive_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a20_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk0_input_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_nios2_oci:the_nios_mcu_nios_cpu_cpu_nios2_oci|nios_mcu_nios_cpu_cpu_nios2_ocimem:the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram_module:nios_mcu_nios_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.operation_mode = "single_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 8;
defparam ram_block1a20.port_a_byte_enable_mask_width = 1;
defparam ram_block1a20.port_a_byte_size = 1;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 255;
defparam ram_block1a20.port_a_logical_ram_depth = 256;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.ram_block_type = "auto";

cycloneive_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a27_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk0_input_clock_enable = "ena0";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_nios2_oci:the_nios_mcu_nios_cpu_cpu_nios2_oci|nios_mcu_nios_cpu_cpu_nios2_ocimem:the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram_module:nios_mcu_nios_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.operation_mode = "single_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 8;
defparam ram_block1a27.port_a_byte_enable_mask_width = 1;
defparam ram_block1a27.port_a_byte_size = 1;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 255;
defparam ram_block1a27.port_a_logical_ram_depth = 256;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.ram_block_type = "auto";

cycloneive_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a28_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.clk0_input_clock_enable = "ena0";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_nios2_oci:the_nios_mcu_nios_cpu_cpu_nios2_oci|nios_mcu_nios_cpu_cpu_nios2_ocimem:the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram_module:nios_mcu_nios_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.operation_mode = "single_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 8;
defparam ram_block1a28.port_a_byte_enable_mask_width = 1;
defparam ram_block1a28.port_a_byte_size = 1;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 255;
defparam ram_block1a28.port_a_logical_ram_depth = 256;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.ram_block_type = "auto";

cycloneive_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a29_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.clk0_input_clock_enable = "ena0";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_nios2_oci:the_nios_mcu_nios_cpu_cpu_nios2_oci|nios_mcu_nios_cpu_cpu_nios2_ocimem:the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram_module:nios_mcu_nios_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.operation_mode = "single_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 8;
defparam ram_block1a29.port_a_byte_enable_mask_width = 1;
defparam ram_block1a29.port_a_byte_size = 1;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 255;
defparam ram_block1a29.port_a_logical_ram_depth = 256;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.ram_block_type = "auto";

cycloneive_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a30_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.clk0_input_clock_enable = "ena0";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_nios2_oci:the_nios_mcu_nios_cpu_cpu_nios2_oci|nios_mcu_nios_cpu_cpu_nios2_ocimem:the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram_module:nios_mcu_nios_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.operation_mode = "single_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 8;
defparam ram_block1a30.port_a_byte_enable_mask_width = 1;
defparam ram_block1a30.port_a_byte_size = 1;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 255;
defparam ram_block1a30.port_a_logical_ram_depth = 256;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.ram_block_type = "auto";

cycloneive_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(!wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a31_PORTADATAOUT_bus),
	.portbdataout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.clk0_input_clock_enable = "ena0";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_nios2_oci:the_nios_mcu_nios_cpu_cpu_nios2_oci|nios_mcu_nios_cpu_cpu_nios2_ocimem:the_nios_mcu_nios_cpu_cpu_nios2_ocimem|nios_mcu_nios_cpu_cpu_ociram_sp_ram_module:nios_mcu_nios_cpu_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_ac71:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.operation_mode = "single_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 8;
defparam ram_block1a31.port_a_byte_enable_mask_width = 1;
defparam ram_block1a31.port_a_byte_size = 1;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 255;
defparam ram_block1a31.port_a_logical_ram_depth = 256;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.ram_block_type = "auto";

endmodule

module nios_mcu_nios_mcu_nios_cpu_cpu_register_bank_a_module (
	q_b_12,
	q_b_11,
	q_b_10,
	q_b_9,
	q_b_8,
	q_b_7,
	q_b_6,
	q_b_5,
	q_b_4,
	q_b_3,
	q_b_2,
	q_b_1,
	q_b_0,
	q_b_15,
	q_b_14,
	q_b_13,
	q_b_31,
	q_b_16,
	q_b_30,
	q_b_29,
	q_b_28,
	q_b_27,
	q_b_26,
	q_b_25,
	q_b_24,
	q_b_23,
	q_b_22,
	q_b_21,
	q_b_20,
	q_b_19,
	q_b_18,
	q_b_17,
	W_rf_wren,
	W_rf_wr_data_0,
	R_dst_regnum_0,
	R_dst_regnum_1,
	R_dst_regnum_2,
	R_dst_regnum_3,
	R_dst_regnum_4,
	W_rf_wr_data_1,
	W_rf_wr_data_2,
	W_rf_wr_data_3,
	W_rf_wr_data_4,
	W_rf_wr_data_5,
	W_rf_wr_data_6,
	W_rf_wr_data_7,
	W_rf_wr_data_12,
	D_iw_27,
	D_iw_28,
	D_iw_29,
	D_iw_30,
	D_iw_31,
	W_rf_wr_data_11,
	W_rf_wr_data_10,
	W_rf_wr_data_9,
	W_rf_wr_data_8,
	W_rf_wr_data_15,
	W_rf_wr_data_14,
	W_rf_wr_data_13,
	W_rf_wr_data_31,
	W_rf_wr_data_16,
	W_rf_wr_data_30,
	W_rf_wr_data_29,
	W_rf_wr_data_28,
	W_rf_wr_data_27,
	W_rf_wr_data_26,
	W_rf_wr_data_25,
	W_rf_wr_data_24,
	W_rf_wr_data_23,
	W_rf_wr_data_22,
	W_rf_wr_data_21,
	W_rf_wr_data_20,
	W_rf_wr_data_19,
	W_rf_wr_data_18,
	W_rf_wr_data_17,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_12;
output 	q_b_11;
output 	q_b_10;
output 	q_b_9;
output 	q_b_8;
output 	q_b_7;
output 	q_b_6;
output 	q_b_5;
output 	q_b_4;
output 	q_b_3;
output 	q_b_2;
output 	q_b_1;
output 	q_b_0;
output 	q_b_15;
output 	q_b_14;
output 	q_b_13;
output 	q_b_31;
output 	q_b_16;
output 	q_b_30;
output 	q_b_29;
output 	q_b_28;
output 	q_b_27;
output 	q_b_26;
output 	q_b_25;
output 	q_b_24;
output 	q_b_23;
output 	q_b_22;
output 	q_b_21;
output 	q_b_20;
output 	q_b_19;
output 	q_b_18;
output 	q_b_17;
input 	W_rf_wren;
input 	W_rf_wr_data_0;
input 	R_dst_regnum_0;
input 	R_dst_regnum_1;
input 	R_dst_regnum_2;
input 	R_dst_regnum_3;
input 	R_dst_regnum_4;
input 	W_rf_wr_data_1;
input 	W_rf_wr_data_2;
input 	W_rf_wr_data_3;
input 	W_rf_wr_data_4;
input 	W_rf_wr_data_5;
input 	W_rf_wr_data_6;
input 	W_rf_wr_data_7;
input 	W_rf_wr_data_12;
input 	D_iw_27;
input 	D_iw_28;
input 	D_iw_29;
input 	D_iw_30;
input 	D_iw_31;
input 	W_rf_wr_data_11;
input 	W_rf_wr_data_10;
input 	W_rf_wr_data_9;
input 	W_rf_wr_data_8;
input 	W_rf_wr_data_15;
input 	W_rf_wr_data_14;
input 	W_rf_wr_data_13;
input 	W_rf_wr_data_31;
input 	W_rf_wr_data_16;
input 	W_rf_wr_data_30;
input 	W_rf_wr_data_29;
input 	W_rf_wr_data_28;
input 	W_rf_wr_data_27;
input 	W_rf_wr_data_26;
input 	W_rf_wr_data_25;
input 	W_rf_wr_data_24;
input 	W_rf_wr_data_23;
input 	W_rf_wr_data_22;
input 	W_rf_wr_data_21;
input 	W_rf_wr_data_20;
input 	W_rf_wr_data_19;
input 	W_rf_wr_data_18;
input 	W_rf_wr_data_17;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nios_mcu_altsyncram_2 the_altsyncram(
	.q_b({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.wren_a(W_rf_wren),
	.data_a({W_rf_wr_data_31,W_rf_wr_data_30,W_rf_wr_data_29,W_rf_wr_data_28,W_rf_wr_data_27,W_rf_wr_data_26,W_rf_wr_data_25,W_rf_wr_data_24,W_rf_wr_data_23,W_rf_wr_data_22,W_rf_wr_data_21,W_rf_wr_data_20,W_rf_wr_data_19,W_rf_wr_data_18,W_rf_wr_data_17,W_rf_wr_data_16,W_rf_wr_data_15,
W_rf_wr_data_14,W_rf_wr_data_13,W_rf_wr_data_12,W_rf_wr_data_11,W_rf_wr_data_10,W_rf_wr_data_9,W_rf_wr_data_8,W_rf_wr_data_7,W_rf_wr_data_6,W_rf_wr_data_5,W_rf_wr_data_4,W_rf_wr_data_3,W_rf_wr_data_2,W_rf_wr_data_1,W_rf_wr_data_0}),
	.address_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,R_dst_regnum_4,R_dst_regnum_3,R_dst_regnum_2,R_dst_regnum_1,R_dst_regnum_0}),
	.address_b({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,D_iw_31,D_iw_30,D_iw_29,D_iw_28,D_iw_27}),
	.clock0(clk_clk));

endmodule

module nios_mcu_altsyncram_2 (
	q_b,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	wren_a;
input 	[31:0] data_a;
input 	[12:0] address_a;
input 	[12:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nios_mcu_altsyncram_6mc1 auto_generated(
	.q_b({q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.wren_a(wren_a),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clock0(clock0));

endmodule

module nios_mcu_altsyncram_6mc1 (
	q_b,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	wren_a;
input 	[31:0] data_a;
input 	[4:0] address_a;
input 	[4:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_a_module:nios_mcu_nios_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_a_module:nios_mcu_nios_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_a_module:nios_mcu_nios_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_a_module:nios_mcu_nios_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_a_module:nios_mcu_nios_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_a_module:nios_mcu_nios_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_a_module:nios_mcu_nios_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_a_module:nios_mcu_nios_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_a_module:nios_mcu_nios_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 5;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 31;
defparam ram_block1a4.port_a_logical_ram_depth = 32;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 5;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 31;
defparam ram_block1a4.port_b_logical_ram_depth = 32;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cycloneive_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_a_module:nios_mcu_nios_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 5;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 31;
defparam ram_block1a3.port_a_logical_ram_depth = 32;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 5;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 31;
defparam ram_block1a3.port_b_logical_ram_depth = 32;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cycloneive_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_a_module:nios_mcu_nios_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 5;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 31;
defparam ram_block1a2.port_a_logical_ram_depth = 32;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 5;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 31;
defparam ram_block1a2.port_b_logical_ram_depth = 32;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cycloneive_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_a_module:nios_mcu_nios_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 5;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 31;
defparam ram_block1a1.port_a_logical_ram_depth = 32;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 5;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 31;
defparam ram_block1a1.port_b_logical_ram_depth = 32;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cycloneive_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_a_module:nios_mcu_nios_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 5;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 31;
defparam ram_block1a0.port_a_logical_ram_depth = 32;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 5;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 31;
defparam ram_block1a0.port_b_logical_ram_depth = 32;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_a_module:nios_mcu_nios_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_a_module:nios_mcu_nios_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_a_module:nios_mcu_nios_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus));
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_a_module:nios_mcu_nios_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 5;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 31;
defparam ram_block1a31.port_a_logical_ram_depth = 32;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock0";
defparam ram_block1a31.port_b_address_width = 5;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 31;
defparam ram_block1a31.port_b_logical_ram_depth = 32;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock0";
defparam ram_block1a31.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_a_module:nios_mcu_nios_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock0";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock0";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus));
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_a_module:nios_mcu_nios_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 5;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 31;
defparam ram_block1a30.port_a_logical_ram_depth = 32;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock0";
defparam ram_block1a30.port_b_address_width = 5;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 31;
defparam ram_block1a30.port_b_logical_ram_depth = 32;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock0";
defparam ram_block1a30.ram_block_type = "auto";

cycloneive_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus));
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_a_module:nios_mcu_nios_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 5;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 31;
defparam ram_block1a29.port_a_logical_ram_depth = 32;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock0";
defparam ram_block1a29.port_b_address_width = 5;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 31;
defparam ram_block1a29.port_b_logical_ram_depth = 32;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock0";
defparam ram_block1a29.ram_block_type = "auto";

cycloneive_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus));
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_a_module:nios_mcu_nios_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 5;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 31;
defparam ram_block1a28.port_a_logical_ram_depth = 32;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock0";
defparam ram_block1a28.port_b_address_width = 5;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 31;
defparam ram_block1a28.port_b_logical_ram_depth = 32;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock0";
defparam ram_block1a28.ram_block_type = "auto";

cycloneive_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus));
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_a_module:nios_mcu_nios_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 5;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 31;
defparam ram_block1a27.port_a_logical_ram_depth = 32;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock0";
defparam ram_block1a27.port_b_address_width = 5;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 31;
defparam ram_block1a27.port_b_logical_ram_depth = 32;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock0";
defparam ram_block1a27.ram_block_type = "auto";

cycloneive_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus));
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_a_module:nios_mcu_nios_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 5;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 31;
defparam ram_block1a26.port_a_logical_ram_depth = 32;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock0";
defparam ram_block1a26.port_b_address_width = 5;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 31;
defparam ram_block1a26.port_b_logical_ram_depth = 32;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock0";
defparam ram_block1a26.ram_block_type = "auto";

cycloneive_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus));
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_a_module:nios_mcu_nios_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 5;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 31;
defparam ram_block1a25.port_a_logical_ram_depth = 32;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock0";
defparam ram_block1a25.port_b_address_width = 5;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 31;
defparam ram_block1a25.port_b_logical_ram_depth = 32;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock0";
defparam ram_block1a25.ram_block_type = "auto";

cycloneive_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus));
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_a_module:nios_mcu_nios_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 5;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 31;
defparam ram_block1a24.port_a_logical_ram_depth = 32;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock0";
defparam ram_block1a24.port_b_address_width = 5;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 31;
defparam ram_block1a24.port_b_logical_ram_depth = 32;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock0";
defparam ram_block1a24.ram_block_type = "auto";

cycloneive_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus));
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_a_module:nios_mcu_nios_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 5;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 31;
defparam ram_block1a23.port_a_logical_ram_depth = 32;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock0";
defparam ram_block1a23.port_b_address_width = 5;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 31;
defparam ram_block1a23.port_b_logical_ram_depth = 32;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock0";
defparam ram_block1a23.ram_block_type = "auto";

cycloneive_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus));
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_a_module:nios_mcu_nios_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 5;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 31;
defparam ram_block1a22.port_a_logical_ram_depth = 32;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock0";
defparam ram_block1a22.port_b_address_width = 5;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 31;
defparam ram_block1a22.port_b_logical_ram_depth = 32;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock0";
defparam ram_block1a22.ram_block_type = "auto";

cycloneive_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus));
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_a_module:nios_mcu_nios_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock0";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock0";
defparam ram_block1a21.ram_block_type = "auto";

cycloneive_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus));
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_a_module:nios_mcu_nios_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock0";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock0";
defparam ram_block1a20.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_a_module:nios_mcu_nios_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock0";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock0";
defparam ram_block1a19.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_a_module:nios_mcu_nios_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock0";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock0";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_a_module:nios_mcu_nios_cpu_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock0";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock0";
defparam ram_block1a17.ram_block_type = "auto";

endmodule

module nios_mcu_nios_mcu_nios_cpu_cpu_register_bank_b_module (
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	q_b_12,
	q_b_11,
	q_b_10,
	q_b_9,
	q_b_8,
	q_b_15,
	q_b_14,
	q_b_13,
	q_b_31,
	q_b_16,
	q_b_30,
	q_b_29,
	q_b_28,
	q_b_27,
	q_b_26,
	q_b_25,
	q_b_24,
	q_b_23,
	q_b_22,
	q_b_21,
	q_b_20,
	q_b_19,
	q_b_18,
	q_b_17,
	W_rf_wren,
	W_rf_wr_data_0,
	R_dst_regnum_0,
	R_dst_regnum_1,
	R_dst_regnum_2,
	R_dst_regnum_3,
	R_dst_regnum_4,
	D_iw_22,
	D_iw_23,
	D_iw_24,
	D_iw_25,
	D_iw_26,
	W_rf_wr_data_1,
	W_rf_wr_data_2,
	W_rf_wr_data_3,
	W_rf_wr_data_4,
	W_rf_wr_data_5,
	W_rf_wr_data_6,
	W_rf_wr_data_7,
	W_rf_wr_data_12,
	W_rf_wr_data_11,
	W_rf_wr_data_10,
	W_rf_wr_data_9,
	W_rf_wr_data_8,
	W_rf_wr_data_15,
	W_rf_wr_data_14,
	W_rf_wr_data_13,
	W_rf_wr_data_31,
	W_rf_wr_data_16,
	W_rf_wr_data_30,
	W_rf_wr_data_29,
	W_rf_wr_data_28,
	W_rf_wr_data_27,
	W_rf_wr_data_26,
	W_rf_wr_data_25,
	W_rf_wr_data_24,
	W_rf_wr_data_23,
	W_rf_wr_data_22,
	W_rf_wr_data_21,
	W_rf_wr_data_20,
	W_rf_wr_data_19,
	W_rf_wr_data_18,
	W_rf_wr_data_17,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
output 	q_b_12;
output 	q_b_11;
output 	q_b_10;
output 	q_b_9;
output 	q_b_8;
output 	q_b_15;
output 	q_b_14;
output 	q_b_13;
output 	q_b_31;
output 	q_b_16;
output 	q_b_30;
output 	q_b_29;
output 	q_b_28;
output 	q_b_27;
output 	q_b_26;
output 	q_b_25;
output 	q_b_24;
output 	q_b_23;
output 	q_b_22;
output 	q_b_21;
output 	q_b_20;
output 	q_b_19;
output 	q_b_18;
output 	q_b_17;
input 	W_rf_wren;
input 	W_rf_wr_data_0;
input 	R_dst_regnum_0;
input 	R_dst_regnum_1;
input 	R_dst_regnum_2;
input 	R_dst_regnum_3;
input 	R_dst_regnum_4;
input 	D_iw_22;
input 	D_iw_23;
input 	D_iw_24;
input 	D_iw_25;
input 	D_iw_26;
input 	W_rf_wr_data_1;
input 	W_rf_wr_data_2;
input 	W_rf_wr_data_3;
input 	W_rf_wr_data_4;
input 	W_rf_wr_data_5;
input 	W_rf_wr_data_6;
input 	W_rf_wr_data_7;
input 	W_rf_wr_data_12;
input 	W_rf_wr_data_11;
input 	W_rf_wr_data_10;
input 	W_rf_wr_data_9;
input 	W_rf_wr_data_8;
input 	W_rf_wr_data_15;
input 	W_rf_wr_data_14;
input 	W_rf_wr_data_13;
input 	W_rf_wr_data_31;
input 	W_rf_wr_data_16;
input 	W_rf_wr_data_30;
input 	W_rf_wr_data_29;
input 	W_rf_wr_data_28;
input 	W_rf_wr_data_27;
input 	W_rf_wr_data_26;
input 	W_rf_wr_data_25;
input 	W_rf_wr_data_24;
input 	W_rf_wr_data_23;
input 	W_rf_wr_data_22;
input 	W_rf_wr_data_21;
input 	W_rf_wr_data_20;
input 	W_rf_wr_data_19;
input 	W_rf_wr_data_18;
input 	W_rf_wr_data_17;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nios_mcu_altsyncram_3 the_altsyncram(
	.q_b({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.wren_a(W_rf_wren),
	.data_a({W_rf_wr_data_31,W_rf_wr_data_30,W_rf_wr_data_29,W_rf_wr_data_28,W_rf_wr_data_27,W_rf_wr_data_26,W_rf_wr_data_25,W_rf_wr_data_24,W_rf_wr_data_23,W_rf_wr_data_22,W_rf_wr_data_21,W_rf_wr_data_20,W_rf_wr_data_19,W_rf_wr_data_18,W_rf_wr_data_17,W_rf_wr_data_16,W_rf_wr_data_15,
W_rf_wr_data_14,W_rf_wr_data_13,W_rf_wr_data_12,W_rf_wr_data_11,W_rf_wr_data_10,W_rf_wr_data_9,W_rf_wr_data_8,W_rf_wr_data_7,W_rf_wr_data_6,W_rf_wr_data_5,W_rf_wr_data_4,W_rf_wr_data_3,W_rf_wr_data_2,W_rf_wr_data_1,W_rf_wr_data_0}),
	.address_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,R_dst_regnum_4,R_dst_regnum_3,R_dst_regnum_2,R_dst_regnum_1,R_dst_regnum_0}),
	.address_b({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,D_iw_26,D_iw_25,D_iw_24,D_iw_23,D_iw_22}),
	.clock0(clk_clk));

endmodule

module nios_mcu_altsyncram_3 (
	q_b,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	wren_a;
input 	[31:0] data_a;
input 	[12:0] address_a;
input 	[12:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nios_mcu_altsyncram_6mc1_1 auto_generated(
	.q_b({q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.wren_a(wren_a),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clock0(clock0));

endmodule

module nios_mcu_altsyncram_6mc1_1 (
	q_b,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	wren_a;
input 	[31:0] data_a;
input 	[4:0] address_a;
input 	[4:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_b_module:nios_mcu_nios_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 5;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 31;
defparam ram_block1a0.port_a_logical_ram_depth = 32;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 5;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 31;
defparam ram_block1a0.port_b_logical_ram_depth = 32;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

cycloneive_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_b_module:nios_mcu_nios_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 5;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 31;
defparam ram_block1a1.port_a_logical_ram_depth = 32;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 5;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 31;
defparam ram_block1a1.port_b_logical_ram_depth = 32;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cycloneive_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_b_module:nios_mcu_nios_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 5;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 31;
defparam ram_block1a2.port_a_logical_ram_depth = 32;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 5;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 31;
defparam ram_block1a2.port_b_logical_ram_depth = 32;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cycloneive_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_b_module:nios_mcu_nios_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 5;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 31;
defparam ram_block1a3.port_a_logical_ram_depth = 32;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 5;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 31;
defparam ram_block1a3.port_b_logical_ram_depth = 32;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cycloneive_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_b_module:nios_mcu_nios_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 5;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 31;
defparam ram_block1a4.port_a_logical_ram_depth = 32;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 5;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 31;
defparam ram_block1a4.port_b_logical_ram_depth = 32;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_b_module:nios_mcu_nios_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_b_module:nios_mcu_nios_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_b_module:nios_mcu_nios_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_b_module:nios_mcu_nios_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_b_module:nios_mcu_nios_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_b_module:nios_mcu_nios_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_b_module:nios_mcu_nios_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_b_module:nios_mcu_nios_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_b_module:nios_mcu_nios_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_b_module:nios_mcu_nios_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_b_module:nios_mcu_nios_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus));
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_b_module:nios_mcu_nios_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 5;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 31;
defparam ram_block1a31.port_a_logical_ram_depth = 32;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock0";
defparam ram_block1a31.port_b_address_width = 5;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 31;
defparam ram_block1a31.port_b_logical_ram_depth = 32;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock0";
defparam ram_block1a31.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_b_module:nios_mcu_nios_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock0";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock0";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus));
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_b_module:nios_mcu_nios_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 5;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 31;
defparam ram_block1a30.port_a_logical_ram_depth = 32;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock0";
defparam ram_block1a30.port_b_address_width = 5;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 31;
defparam ram_block1a30.port_b_logical_ram_depth = 32;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock0";
defparam ram_block1a30.ram_block_type = "auto";

cycloneive_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus));
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_b_module:nios_mcu_nios_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 5;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 31;
defparam ram_block1a29.port_a_logical_ram_depth = 32;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock0";
defparam ram_block1a29.port_b_address_width = 5;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 31;
defparam ram_block1a29.port_b_logical_ram_depth = 32;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock0";
defparam ram_block1a29.ram_block_type = "auto";

cycloneive_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus));
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_b_module:nios_mcu_nios_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 5;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 31;
defparam ram_block1a28.port_a_logical_ram_depth = 32;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock0";
defparam ram_block1a28.port_b_address_width = 5;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 31;
defparam ram_block1a28.port_b_logical_ram_depth = 32;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock0";
defparam ram_block1a28.ram_block_type = "auto";

cycloneive_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus));
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_b_module:nios_mcu_nios_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 5;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 31;
defparam ram_block1a27.port_a_logical_ram_depth = 32;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock0";
defparam ram_block1a27.port_b_address_width = 5;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 31;
defparam ram_block1a27.port_b_logical_ram_depth = 32;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock0";
defparam ram_block1a27.ram_block_type = "auto";

cycloneive_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus));
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_b_module:nios_mcu_nios_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 5;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 31;
defparam ram_block1a26.port_a_logical_ram_depth = 32;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock0";
defparam ram_block1a26.port_b_address_width = 5;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 31;
defparam ram_block1a26.port_b_logical_ram_depth = 32;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock0";
defparam ram_block1a26.ram_block_type = "auto";

cycloneive_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus));
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_b_module:nios_mcu_nios_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 5;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 31;
defparam ram_block1a25.port_a_logical_ram_depth = 32;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock0";
defparam ram_block1a25.port_b_address_width = 5;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 31;
defparam ram_block1a25.port_b_logical_ram_depth = 32;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock0";
defparam ram_block1a25.ram_block_type = "auto";

cycloneive_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus));
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_b_module:nios_mcu_nios_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 5;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 31;
defparam ram_block1a24.port_a_logical_ram_depth = 32;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock0";
defparam ram_block1a24.port_b_address_width = 5;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 31;
defparam ram_block1a24.port_b_logical_ram_depth = 32;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock0";
defparam ram_block1a24.ram_block_type = "auto";

cycloneive_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus));
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_b_module:nios_mcu_nios_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 5;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 31;
defparam ram_block1a23.port_a_logical_ram_depth = 32;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock0";
defparam ram_block1a23.port_b_address_width = 5;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 31;
defparam ram_block1a23.port_b_logical_ram_depth = 32;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock0";
defparam ram_block1a23.ram_block_type = "auto";

cycloneive_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus));
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_b_module:nios_mcu_nios_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 5;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 31;
defparam ram_block1a22.port_a_logical_ram_depth = 32;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock0";
defparam ram_block1a22.port_b_address_width = 5;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 31;
defparam ram_block1a22.port_b_logical_ram_depth = 32;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock0";
defparam ram_block1a22.ram_block_type = "auto";

cycloneive_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus));
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_b_module:nios_mcu_nios_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock0";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock0";
defparam ram_block1a21.ram_block_type = "auto";

cycloneive_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus));
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_b_module:nios_mcu_nios_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock0";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock0";
defparam ram_block1a20.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_b_module:nios_mcu_nios_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock0";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock0";
defparam ram_block1a19.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_b_module:nios_mcu_nios_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock0";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock0";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "nios_mcu_nios_cpu:nios_cpu|nios_mcu_nios_cpu_cpu:cpu|nios_mcu_nios_cpu_cpu_register_bank_b_module:nios_mcu_nios_cpu_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_6mc1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock0";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock0";
defparam ram_block1a17.ram_block_type = "auto";

endmodule

module nios_mcu_nios_mcu_onchip_ram (
	W_alu_result_12,
	W_alu_result_14,
	W_alu_result_13,
	W_alu_result_11,
	W_alu_result_10,
	W_alu_result_9,
	W_alu_result_8,
	W_alu_result_7,
	W_alu_result_6,
	W_alu_result_5,
	W_alu_result_4,
	W_alu_result_3,
	W_alu_result_2,
	q_a_0,
	q_b_0,
	q_a_22,
	q_b_22,
	q_a_23,
	q_b_23,
	q_a_24,
	q_b_24,
	q_a_25,
	q_b_25,
	q_a_26,
	q_b_26,
	q_a_11,
	q_b_11,
	q_a_13,
	q_b_13,
	q_a_16,
	q_b_16,
	q_a_12,
	q_b_12,
	q_a_1,
	q_b_1,
	q_a_3,
	q_b_3,
	q_a_2,
	q_b_2,
	q_a_5,
	q_b_5,
	q_a_4,
	q_b_4,
	q_a_14,
	q_b_14,
	q_a_15,
	q_b_15,
	q_a_18,
	q_b_18,
	q_a_17,
	q_b_17,
	q_a_10,
	q_b_10,
	q_a_9,
	q_b_9,
	q_a_8,
	q_b_8,
	q_a_7,
	q_b_7,
	q_a_6,
	q_b_6,
	q_a_21,
	q_b_21,
	q_a_19,
	q_b_19,
	q_a_20,
	q_b_20,
	d_writedata_24,
	d_writedata_25,
	d_writedata_26,
	q_a_27,
	q_b_27,
	q_a_28,
	q_b_28,
	q_a_29,
	q_b_29,
	q_a_30,
	q_b_30,
	q_a_31,
	q_b_31,
	d_writedata_27,
	d_writedata_28,
	d_writedata_29,
	d_writedata_30,
	d_writedata_31,
	d_writedata_0,
	rst1,
	d_writedata_1,
	d_writedata_2,
	d_writedata_3,
	d_writedata_4,
	d_writedata_5,
	d_writedata_6,
	d_writedata_7,
	m0_write,
	src_channel_4,
	mem_used_1,
	F_pc_10,
	F_pc_9,
	F_pc_8,
	F_pc_7,
	F_pc_6,
	F_pc_5,
	F_pc_4,
	F_pc_3,
	F_pc_2,
	F_pc_1,
	F_pc_0,
	F_pc_12,
	F_pc_11,
	r_early_rst,
	d_byteenable_0,
	d_writedata_22,
	d_byteenable_2,
	d_writedata_23,
	d_byteenable_3,
	d_writedata_11,
	d_byteenable_1,
	d_writedata_13,
	d_writedata_16,
	d_writedata_12,
	d_writedata_14,
	d_writedata_15,
	d_writedata_18,
	d_writedata_17,
	d_writedata_10,
	d_writedata_9,
	d_writedata_8,
	d_writedata_21,
	d_writedata_19,
	d_writedata_20,
	GND_port,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_12;
input 	W_alu_result_14;
input 	W_alu_result_13;
input 	W_alu_result_11;
input 	W_alu_result_10;
input 	W_alu_result_9;
input 	W_alu_result_8;
input 	W_alu_result_7;
input 	W_alu_result_6;
input 	W_alu_result_5;
input 	W_alu_result_4;
input 	W_alu_result_3;
input 	W_alu_result_2;
output 	q_a_0;
output 	q_b_0;
output 	q_a_22;
output 	q_b_22;
output 	q_a_23;
output 	q_b_23;
output 	q_a_24;
output 	q_b_24;
output 	q_a_25;
output 	q_b_25;
output 	q_a_26;
output 	q_b_26;
output 	q_a_11;
output 	q_b_11;
output 	q_a_13;
output 	q_b_13;
output 	q_a_16;
output 	q_b_16;
output 	q_a_12;
output 	q_b_12;
output 	q_a_1;
output 	q_b_1;
output 	q_a_3;
output 	q_b_3;
output 	q_a_2;
output 	q_b_2;
output 	q_a_5;
output 	q_b_5;
output 	q_a_4;
output 	q_b_4;
output 	q_a_14;
output 	q_b_14;
output 	q_a_15;
output 	q_b_15;
output 	q_a_18;
output 	q_b_18;
output 	q_a_17;
output 	q_b_17;
output 	q_a_10;
output 	q_b_10;
output 	q_a_9;
output 	q_b_9;
output 	q_a_8;
output 	q_b_8;
output 	q_a_7;
output 	q_b_7;
output 	q_a_6;
output 	q_b_6;
output 	q_a_21;
output 	q_b_21;
output 	q_a_19;
output 	q_b_19;
output 	q_a_20;
output 	q_b_20;
input 	d_writedata_24;
input 	d_writedata_25;
input 	d_writedata_26;
output 	q_a_27;
output 	q_b_27;
output 	q_a_28;
output 	q_b_28;
output 	q_a_29;
output 	q_b_29;
output 	q_a_30;
output 	q_b_30;
output 	q_a_31;
output 	q_b_31;
input 	d_writedata_27;
input 	d_writedata_28;
input 	d_writedata_29;
input 	d_writedata_30;
input 	d_writedata_31;
input 	d_writedata_0;
input 	rst1;
input 	d_writedata_1;
input 	d_writedata_2;
input 	d_writedata_3;
input 	d_writedata_4;
input 	d_writedata_5;
input 	d_writedata_6;
input 	d_writedata_7;
input 	m0_write;
input 	src_channel_4;
input 	mem_used_1;
input 	F_pc_10;
input 	F_pc_9;
input 	F_pc_8;
input 	F_pc_7;
input 	F_pc_6;
input 	F_pc_5;
input 	F_pc_4;
input 	F_pc_3;
input 	F_pc_2;
input 	F_pc_1;
input 	F_pc_0;
input 	F_pc_12;
input 	F_pc_11;
input 	r_early_rst;
input 	d_byteenable_0;
input 	d_writedata_22;
input 	d_byteenable_2;
input 	d_writedata_23;
input 	d_byteenable_3;
input 	d_writedata_11;
input 	d_byteenable_1;
input 	d_writedata_13;
input 	d_writedata_16;
input 	d_writedata_12;
input 	d_writedata_14;
input 	d_writedata_15;
input 	d_writedata_18;
input 	d_writedata_17;
input 	d_writedata_10;
input 	d_writedata_9;
input 	d_writedata_8;
input 	d_writedata_21;
input 	d_writedata_19;
input 	d_writedata_20;
input 	GND_port;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wren2~0_combout ;


nios_mcu_altsyncram_4 the_altsyncram(
	.address_b({W_alu_result_14,W_alu_result_13,W_alu_result_12,W_alu_result_11,W_alu_result_10,W_alu_result_9,W_alu_result_8,W_alu_result_7,W_alu_result_6,W_alu_result_5,W_alu_result_4,W_alu_result_3,W_alu_result_2}),
	.q_a({q_a_31,q_a_30,q_a_29,q_a_28,q_a_27,q_a_26,q_a_25,q_a_24,q_a_23,q_a_22,q_a_21,q_a_20,q_a_19,q_a_18,q_a_17,q_a_16,q_a_15,q_a_14,q_a_13,q_a_12,q_a_11,q_a_10,q_a_9,q_a_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.q_b({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.data_b({d_writedata_31,d_writedata_30,d_writedata_29,d_writedata_28,d_writedata_27,d_writedata_26,d_writedata_25,d_writedata_24,d_writedata_23,d_writedata_22,d_writedata_21,d_writedata_20,d_writedata_19,d_writedata_18,d_writedata_17,d_writedata_16,d_writedata_15,d_writedata_14,
d_writedata_13,d_writedata_12,d_writedata_11,d_writedata_10,d_writedata_9,d_writedata_8,d_writedata_7,d_writedata_6,d_writedata_5,d_writedata_4,d_writedata_3,d_writedata_2,d_writedata_1,d_writedata_0}),
	.address_a({F_pc_12,F_pc_11,F_pc_10,F_pc_9,F_pc_8,F_pc_7,F_pc_6,F_pc_5,F_pc_4,F_pc_3,F_pc_2,F_pc_1,F_pc_0}),
	.clocken0(r_early_rst),
	.wren_b(\wren2~0_combout ),
	.byteena_b({d_byteenable_3,d_byteenable_2,d_byteenable_1,d_byteenable_0}),
	.data_a({GND_port,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.clock0(clk_clk));

cycloneive_lcell_comb \wren2~0 (
	.dataa(mem_used_1),
	.datab(rst1),
	.datac(m0_write),
	.datad(src_channel_4),
	.cin(gnd),
	.combout(\wren2~0_combout ),
	.cout());
defparam \wren2~0 .lut_mask = 16'hFFFD;
defparam \wren2~0 .sum_lutc_input = "datac";

endmodule

module nios_mcu_altsyncram_4 (
	address_b,
	q_a,
	q_b,
	data_b,
	address_a,
	clocken0,
	wren_b,
	byteena_b,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
input 	[12:0] address_b;
output 	[31:0] q_a;
output 	[31:0] q_b;
input 	[31:0] data_b;
input 	[12:0] address_a;
input 	clocken0;
input 	wren_b;
input 	[3:0] byteena_b;
input 	[31:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nios_mcu_altsyncram_h232 auto_generated(
	.address_b({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.q_a({q_a[31],q_a[30],q_a[29],q_a[28],q_a[27],q_a[26],q_a[25],q_a[24],q_a[23],q_a[22],q_a[21],q_a[20],q_a[19],q_a[18],q_a[17],q_a[16],q_a[15],q_a[14],q_a[13],q_a[12],q_a[11],q_a[10],q_a[9],q_a[8],q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.q_b({q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.data_b({data_b[31],data_b[30],data_b[29],data_b[28],data_b[27],data_b[26],data_b[25],data_b[24],data_b[23],data_b[22],data_b[21],data_b[20],data_b[19],data_b[18],data_b[17],data_b[16],data_b[15],data_b[14],data_b[13],data_b[12],data_b[11],data_b[10],data_b[9],data_b[8],data_b[7],data_b[6],data_b[5],data_b[4],data_b[3],data_b[2],data_b[1],data_b[0]}),
	.address_a({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.clocken0(clocken0),
	.wren_b(wren_b),
	.byteena_b({byteena_b[3],byteena_b[2],byteena_b[1],byteena_b[0]}),
	.data_a({data_a[31],data_a[31],data_a[31],data_a[31],data_a[31],data_a[31],data_a[31],data_a[31],data_a[31],data_a[31],data_a[31],data_a[31],data_a[31],data_a[31],data_a[31],data_a[31],data_a[31],data_a[31],data_a[31],data_a[31],data_a[31],data_a[31],data_a[31],data_a[31],data_a[31],data_a[31],data_a[31],data_a[31],data_a[31],data_a[31],data_a[31],data_a[31]}),
	.clock0(clock0));

endmodule

module nios_mcu_altsyncram_h232 (
	address_b,
	q_a,
	q_b,
	data_b,
	address_a,
	clocken0,
	wren_b,
	byteena_b,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
input 	[12:0] address_b;
output 	[31:0] q_a;
output 	[31:0] q_b;
input 	[31:0] data_b;
input 	[12:0] address_a;
input 	clocken0;
input 	wren_b;
input 	[3:0] byteena_b;
input 	[31:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTADATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTADATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTADATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTADATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTADATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTADATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTADATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTADATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTADATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTADATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTADATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTADATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTADATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTADATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTADATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTADATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTADATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTADATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTADATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTADATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTADATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTADATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_a[22] = ram_block1a22_PORTADATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_a[23] = ram_block1a23_PORTADATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_a[24] = ram_block1a24_PORTADATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_a[25] = ram_block1a25_PORTADATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_a[26] = ram_block1a26_PORTADATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_a[11] = ram_block1a11_PORTADATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_a[13] = ram_block1a13_PORTADATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_a[16] = ram_block1a16_PORTADATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_a[12] = ram_block1a12_PORTADATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_a[14] = ram_block1a14_PORTADATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_a[15] = ram_block1a15_PORTADATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_a[18] = ram_block1a18_PORTADATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_a[17] = ram_block1a17_PORTADATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_a[10] = ram_block1a10_PORTADATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_a[9] = ram_block1a9_PORTADATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_a[8] = ram_block1a8_PORTADATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_a[21] = ram_block1a21_PORTADATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_a[19] = ram_block1a19_PORTADATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_a[20] = ram_block1a20_PORTADATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_a[27] = ram_block1a27_PORTADATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_a[28] = ram_block1a28_PORTADATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_a[29] = ram_block1a29_PORTADATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_a[30] = ram_block1a30_PORTADATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_a[31] = ram_block1a31_PORTADATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a0(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[0]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "nios_mcu_onchip_ram.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "nios_mcu_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_h232:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "bidir_dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 13;
defparam ram_block1a0.port_a_byte_enable_mask_width = 1;
defparam ram_block1a0.port_a_byte_size = 1;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 8191;
defparam ram_block1a0.port_a_logical_ram_depth = 8192;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 13;
defparam ram_block1a0.port_b_byte_enable_clock = "clock0";
defparam ram_block1a0.port_b_byte_enable_mask_width = 1;
defparam ram_block1a0.port_b_byte_size = 1;
defparam ram_block1a0.port_b_data_in_clock = "clock0";
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 8191;
defparam ram_block1a0.port_b_logical_ram_depth = 8192;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.port_b_write_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a0.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a0.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a0.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneive_ram_block ram_block1a22(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[22]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a22_PORTADATAOUT_bus),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus));
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk0_input_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.init_file = "nios_mcu_onchip_ram.hex";
defparam ram_block1a22.init_file_layout = "port_a";
defparam ram_block1a22.logical_ram_name = "nios_mcu_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_h232:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "bidir_dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 13;
defparam ram_block1a22.port_a_byte_enable_mask_width = 1;
defparam ram_block1a22.port_a_byte_size = 1;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 8191;
defparam ram_block1a22.port_a_logical_ram_depth = 8192;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock0";
defparam ram_block1a22.port_b_address_width = 13;
defparam ram_block1a22.port_b_byte_enable_clock = "clock0";
defparam ram_block1a22.port_b_byte_enable_mask_width = 1;
defparam ram_block1a22.port_b_byte_size = 1;
defparam ram_block1a22.port_b_data_in_clock = "clock0";
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 8191;
defparam ram_block1a22.port_b_logical_ram_depth = 8192;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock0";
defparam ram_block1a22.port_b_write_enable_clock = "clock0";
defparam ram_block1a22.ram_block_type = "auto";
defparam ram_block1a22.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a22.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a22.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a22.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneive_ram_block ram_block1a23(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[23]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a23_PORTADATAOUT_bus),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus));
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk0_input_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.init_file = "nios_mcu_onchip_ram.hex";
defparam ram_block1a23.init_file_layout = "port_a";
defparam ram_block1a23.logical_ram_name = "nios_mcu_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_h232:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "bidir_dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 13;
defparam ram_block1a23.port_a_byte_enable_mask_width = 1;
defparam ram_block1a23.port_a_byte_size = 1;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 8191;
defparam ram_block1a23.port_a_logical_ram_depth = 8192;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock0";
defparam ram_block1a23.port_b_address_width = 13;
defparam ram_block1a23.port_b_byte_enable_clock = "clock0";
defparam ram_block1a23.port_b_byte_enable_mask_width = 1;
defparam ram_block1a23.port_b_byte_size = 1;
defparam ram_block1a23.port_b_data_in_clock = "clock0";
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 8191;
defparam ram_block1a23.port_b_logical_ram_depth = 8192;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock0";
defparam ram_block1a23.port_b_write_enable_clock = "clock0";
defparam ram_block1a23.ram_block_type = "auto";
defparam ram_block1a23.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a23.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a23.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a23.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneive_ram_block ram_block1a24(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[24]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a24_PORTADATAOUT_bus),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus));
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk0_input_clock_enable = "ena0";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.init_file = "nios_mcu_onchip_ram.hex";
defparam ram_block1a24.init_file_layout = "port_a";
defparam ram_block1a24.logical_ram_name = "nios_mcu_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_h232:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "bidir_dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 13;
defparam ram_block1a24.port_a_byte_enable_mask_width = 1;
defparam ram_block1a24.port_a_byte_size = 1;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 8191;
defparam ram_block1a24.port_a_logical_ram_depth = 8192;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock0";
defparam ram_block1a24.port_b_address_width = 13;
defparam ram_block1a24.port_b_byte_enable_clock = "clock0";
defparam ram_block1a24.port_b_byte_enable_mask_width = 1;
defparam ram_block1a24.port_b_byte_size = 1;
defparam ram_block1a24.port_b_data_in_clock = "clock0";
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 8191;
defparam ram_block1a24.port_b_logical_ram_depth = 8192;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock0";
defparam ram_block1a24.port_b_write_enable_clock = "clock0";
defparam ram_block1a24.ram_block_type = "auto";
defparam ram_block1a24.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a24.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a24.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a24.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneive_ram_block ram_block1a25(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[25]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a25_PORTADATAOUT_bus),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus));
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk0_input_clock_enable = "ena0";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.init_file = "nios_mcu_onchip_ram.hex";
defparam ram_block1a25.init_file_layout = "port_a";
defparam ram_block1a25.logical_ram_name = "nios_mcu_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_h232:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "bidir_dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 13;
defparam ram_block1a25.port_a_byte_enable_mask_width = 1;
defparam ram_block1a25.port_a_byte_size = 1;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 8191;
defparam ram_block1a25.port_a_logical_ram_depth = 8192;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock0";
defparam ram_block1a25.port_b_address_width = 13;
defparam ram_block1a25.port_b_byte_enable_clock = "clock0";
defparam ram_block1a25.port_b_byte_enable_mask_width = 1;
defparam ram_block1a25.port_b_byte_size = 1;
defparam ram_block1a25.port_b_data_in_clock = "clock0";
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 8191;
defparam ram_block1a25.port_b_logical_ram_depth = 8192;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock0";
defparam ram_block1a25.port_b_write_enable_clock = "clock0";
defparam ram_block1a25.ram_block_type = "auto";
defparam ram_block1a25.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a25.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a25.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a25.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneive_ram_block ram_block1a26(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[26]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a26_PORTADATAOUT_bus),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus));
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk0_input_clock_enable = "ena0";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.init_file = "nios_mcu_onchip_ram.hex";
defparam ram_block1a26.init_file_layout = "port_a";
defparam ram_block1a26.logical_ram_name = "nios_mcu_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_h232:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "bidir_dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 13;
defparam ram_block1a26.port_a_byte_enable_mask_width = 1;
defparam ram_block1a26.port_a_byte_size = 1;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 8191;
defparam ram_block1a26.port_a_logical_ram_depth = 8192;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock0";
defparam ram_block1a26.port_b_address_width = 13;
defparam ram_block1a26.port_b_byte_enable_clock = "clock0";
defparam ram_block1a26.port_b_byte_enable_mask_width = 1;
defparam ram_block1a26.port_b_byte_size = 1;
defparam ram_block1a26.port_b_data_in_clock = "clock0";
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 8191;
defparam ram_block1a26.port_b_logical_ram_depth = 8192;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock0";
defparam ram_block1a26.port_b_write_enable_clock = "clock0";
defparam ram_block1a26.ram_block_type = "auto";
defparam ram_block1a26.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a26.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a26.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a26.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneive_ram_block ram_block1a11(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[11]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a11_PORTADATAOUT_bus),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.init_file = "nios_mcu_onchip_ram.hex";
defparam ram_block1a11.init_file_layout = "port_a";
defparam ram_block1a11.logical_ram_name = "nios_mcu_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_h232:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "bidir_dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 13;
defparam ram_block1a11.port_a_byte_enable_mask_width = 1;
defparam ram_block1a11.port_a_byte_size = 1;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 8191;
defparam ram_block1a11.port_a_logical_ram_depth = 8192;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 13;
defparam ram_block1a11.port_b_byte_enable_clock = "clock0";
defparam ram_block1a11.port_b_byte_enable_mask_width = 1;
defparam ram_block1a11.port_b_byte_size = 1;
defparam ram_block1a11.port_b_data_in_clock = "clock0";
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 8191;
defparam ram_block1a11.port_b_logical_ram_depth = 8192;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.port_b_write_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";
defparam ram_block1a11.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a11.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a11.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a11.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneive_ram_block ram_block1a13(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[13]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a13_PORTADATAOUT_bus),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.init_file = "nios_mcu_onchip_ram.hex";
defparam ram_block1a13.init_file_layout = "port_a";
defparam ram_block1a13.logical_ram_name = "nios_mcu_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_h232:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "bidir_dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 13;
defparam ram_block1a13.port_a_byte_enable_mask_width = 1;
defparam ram_block1a13.port_a_byte_size = 1;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 8191;
defparam ram_block1a13.port_a_logical_ram_depth = 8192;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 13;
defparam ram_block1a13.port_b_byte_enable_clock = "clock0";
defparam ram_block1a13.port_b_byte_enable_mask_width = 1;
defparam ram_block1a13.port_b_byte_size = 1;
defparam ram_block1a13.port_b_data_in_clock = "clock0";
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 8191;
defparam ram_block1a13.port_b_logical_ram_depth = 8192;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.port_b_write_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";
defparam ram_block1a13.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a13.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a13.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a13.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneive_ram_block ram_block1a16(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[16]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a16_PORTADATAOUT_bus),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.init_file = "nios_mcu_onchip_ram.hex";
defparam ram_block1a16.init_file_layout = "port_a";
defparam ram_block1a16.logical_ram_name = "nios_mcu_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_h232:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "bidir_dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 13;
defparam ram_block1a16.port_a_byte_enable_mask_width = 1;
defparam ram_block1a16.port_a_byte_size = 1;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 8191;
defparam ram_block1a16.port_a_logical_ram_depth = 8192;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock0";
defparam ram_block1a16.port_b_address_width = 13;
defparam ram_block1a16.port_b_byte_enable_clock = "clock0";
defparam ram_block1a16.port_b_byte_enable_mask_width = 1;
defparam ram_block1a16.port_b_byte_size = 1;
defparam ram_block1a16.port_b_data_in_clock = "clock0";
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 8191;
defparam ram_block1a16.port_b_logical_ram_depth = 8192;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock0";
defparam ram_block1a16.port_b_write_enable_clock = "clock0";
defparam ram_block1a16.ram_block_type = "auto";
defparam ram_block1a16.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a16.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a16.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a16.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneive_ram_block ram_block1a12(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[12]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a12_PORTADATAOUT_bus),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.init_file = "nios_mcu_onchip_ram.hex";
defparam ram_block1a12.init_file_layout = "port_a";
defparam ram_block1a12.logical_ram_name = "nios_mcu_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_h232:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "bidir_dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 13;
defparam ram_block1a12.port_a_byte_enable_mask_width = 1;
defparam ram_block1a12.port_a_byte_size = 1;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 8191;
defparam ram_block1a12.port_a_logical_ram_depth = 8192;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 13;
defparam ram_block1a12.port_b_byte_enable_clock = "clock0";
defparam ram_block1a12.port_b_byte_enable_mask_width = 1;
defparam ram_block1a12.port_b_byte_size = 1;
defparam ram_block1a12.port_b_data_in_clock = "clock0";
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 8191;
defparam ram_block1a12.port_b_logical_ram_depth = 8192;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.port_b_write_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";
defparam ram_block1a12.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a12.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a12.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a12.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneive_ram_block ram_block1a1(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[1]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "nios_mcu_onchip_ram.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "nios_mcu_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_h232:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "bidir_dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 13;
defparam ram_block1a1.port_a_byte_enable_mask_width = 1;
defparam ram_block1a1.port_a_byte_size = 1;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 8191;
defparam ram_block1a1.port_a_logical_ram_depth = 8192;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 13;
defparam ram_block1a1.port_b_byte_enable_clock = "clock0";
defparam ram_block1a1.port_b_byte_enable_mask_width = 1;
defparam ram_block1a1.port_b_byte_size = 1;
defparam ram_block1a1.port_b_data_in_clock = "clock0";
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 8191;
defparam ram_block1a1.port_b_logical_ram_depth = 8192;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.port_b_write_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a1.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a1.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a1.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneive_ram_block ram_block1a3(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[3]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "nios_mcu_onchip_ram.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "nios_mcu_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_h232:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "bidir_dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 13;
defparam ram_block1a3.port_a_byte_enable_mask_width = 1;
defparam ram_block1a3.port_a_byte_size = 1;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 8191;
defparam ram_block1a3.port_a_logical_ram_depth = 8192;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 13;
defparam ram_block1a3.port_b_byte_enable_clock = "clock0";
defparam ram_block1a3.port_b_byte_enable_mask_width = 1;
defparam ram_block1a3.port_b_byte_size = 1;
defparam ram_block1a3.port_b_data_in_clock = "clock0";
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 8191;
defparam ram_block1a3.port_b_logical_ram_depth = 8192;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.port_b_write_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a3.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a3.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a3.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneive_ram_block ram_block1a2(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[2]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "nios_mcu_onchip_ram.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "nios_mcu_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_h232:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "bidir_dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 13;
defparam ram_block1a2.port_a_byte_enable_mask_width = 1;
defparam ram_block1a2.port_a_byte_size = 1;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 8191;
defparam ram_block1a2.port_a_logical_ram_depth = 8192;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 13;
defparam ram_block1a2.port_b_byte_enable_clock = "clock0";
defparam ram_block1a2.port_b_byte_enable_mask_width = 1;
defparam ram_block1a2.port_b_byte_size = 1;
defparam ram_block1a2.port_b_data_in_clock = "clock0";
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 8191;
defparam ram_block1a2.port_b_logical_ram_depth = 8192;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.port_b_write_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a2.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a2.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a2.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneive_ram_block ram_block1a5(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[5]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "nios_mcu_onchip_ram.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "nios_mcu_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_h232:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "bidir_dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 13;
defparam ram_block1a5.port_a_byte_enable_mask_width = 1;
defparam ram_block1a5.port_a_byte_size = 1;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 8191;
defparam ram_block1a5.port_a_logical_ram_depth = 8192;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 13;
defparam ram_block1a5.port_b_byte_enable_clock = "clock0";
defparam ram_block1a5.port_b_byte_enable_mask_width = 1;
defparam ram_block1a5.port_b_byte_size = 1;
defparam ram_block1a5.port_b_data_in_clock = "clock0";
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 8191;
defparam ram_block1a5.port_b_logical_ram_depth = 8192;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.port_b_write_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a5.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a5.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a5.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneive_ram_block ram_block1a4(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[4]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "nios_mcu_onchip_ram.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "nios_mcu_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_h232:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "bidir_dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 13;
defparam ram_block1a4.port_a_byte_enable_mask_width = 1;
defparam ram_block1a4.port_a_byte_size = 1;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 8191;
defparam ram_block1a4.port_a_logical_ram_depth = 8192;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 13;
defparam ram_block1a4.port_b_byte_enable_clock = "clock0";
defparam ram_block1a4.port_b_byte_enable_mask_width = 1;
defparam ram_block1a4.port_b_byte_size = 1;
defparam ram_block1a4.port_b_data_in_clock = "clock0";
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 8191;
defparam ram_block1a4.port_b_logical_ram_depth = 8192;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.port_b_write_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a4.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a4.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a4.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneive_ram_block ram_block1a14(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[14]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a14_PORTADATAOUT_bus),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.init_file = "nios_mcu_onchip_ram.hex";
defparam ram_block1a14.init_file_layout = "port_a";
defparam ram_block1a14.logical_ram_name = "nios_mcu_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_h232:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "bidir_dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 13;
defparam ram_block1a14.port_a_byte_enable_mask_width = 1;
defparam ram_block1a14.port_a_byte_size = 1;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 8191;
defparam ram_block1a14.port_a_logical_ram_depth = 8192;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 13;
defparam ram_block1a14.port_b_byte_enable_clock = "clock0";
defparam ram_block1a14.port_b_byte_enable_mask_width = 1;
defparam ram_block1a14.port_b_byte_size = 1;
defparam ram_block1a14.port_b_data_in_clock = "clock0";
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 8191;
defparam ram_block1a14.port_b_logical_ram_depth = 8192;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.port_b_write_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";
defparam ram_block1a14.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a14.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a14.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a14.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneive_ram_block ram_block1a15(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[15]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a15_PORTADATAOUT_bus),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.init_file = "nios_mcu_onchip_ram.hex";
defparam ram_block1a15.init_file_layout = "port_a";
defparam ram_block1a15.logical_ram_name = "nios_mcu_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_h232:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "bidir_dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 13;
defparam ram_block1a15.port_a_byte_enable_mask_width = 1;
defparam ram_block1a15.port_a_byte_size = 1;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 8191;
defparam ram_block1a15.port_a_logical_ram_depth = 8192;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 13;
defparam ram_block1a15.port_b_byte_enable_clock = "clock0";
defparam ram_block1a15.port_b_byte_enable_mask_width = 1;
defparam ram_block1a15.port_b_byte_size = 1;
defparam ram_block1a15.port_b_data_in_clock = "clock0";
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 8191;
defparam ram_block1a15.port_b_logical_ram_depth = 8192;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.port_b_write_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";
defparam ram_block1a15.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a15.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a15.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a15.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneive_ram_block ram_block1a18(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[18]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a18_PORTADATAOUT_bus),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.init_file = "nios_mcu_onchip_ram.hex";
defparam ram_block1a18.init_file_layout = "port_a";
defparam ram_block1a18.logical_ram_name = "nios_mcu_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_h232:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "bidir_dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 13;
defparam ram_block1a18.port_a_byte_enable_mask_width = 1;
defparam ram_block1a18.port_a_byte_size = 1;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 8191;
defparam ram_block1a18.port_a_logical_ram_depth = 8192;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock0";
defparam ram_block1a18.port_b_address_width = 13;
defparam ram_block1a18.port_b_byte_enable_clock = "clock0";
defparam ram_block1a18.port_b_byte_enable_mask_width = 1;
defparam ram_block1a18.port_b_byte_size = 1;
defparam ram_block1a18.port_b_data_in_clock = "clock0";
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 8191;
defparam ram_block1a18.port_b_logical_ram_depth = 8192;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock0";
defparam ram_block1a18.port_b_write_enable_clock = "clock0";
defparam ram_block1a18.ram_block_type = "auto";
defparam ram_block1a18.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a18.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a18.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a18.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneive_ram_block ram_block1a17(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[17]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a17_PORTADATAOUT_bus),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.init_file = "nios_mcu_onchip_ram.hex";
defparam ram_block1a17.init_file_layout = "port_a";
defparam ram_block1a17.logical_ram_name = "nios_mcu_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_h232:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "bidir_dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 13;
defparam ram_block1a17.port_a_byte_enable_mask_width = 1;
defparam ram_block1a17.port_a_byte_size = 1;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 8191;
defparam ram_block1a17.port_a_logical_ram_depth = 8192;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock0";
defparam ram_block1a17.port_b_address_width = 13;
defparam ram_block1a17.port_b_byte_enable_clock = "clock0";
defparam ram_block1a17.port_b_byte_enable_mask_width = 1;
defparam ram_block1a17.port_b_byte_size = 1;
defparam ram_block1a17.port_b_data_in_clock = "clock0";
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 8191;
defparam ram_block1a17.port_b_logical_ram_depth = 8192;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock0";
defparam ram_block1a17.port_b_write_enable_clock = "clock0";
defparam ram_block1a17.ram_block_type = "auto";
defparam ram_block1a17.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a17.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a17.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a17.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneive_ram_block ram_block1a10(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[10]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a10_PORTADATAOUT_bus),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.init_file = "nios_mcu_onchip_ram.hex";
defparam ram_block1a10.init_file_layout = "port_a";
defparam ram_block1a10.logical_ram_name = "nios_mcu_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_h232:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "bidir_dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 13;
defparam ram_block1a10.port_a_byte_enable_mask_width = 1;
defparam ram_block1a10.port_a_byte_size = 1;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 8191;
defparam ram_block1a10.port_a_logical_ram_depth = 8192;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 13;
defparam ram_block1a10.port_b_byte_enable_clock = "clock0";
defparam ram_block1a10.port_b_byte_enable_mask_width = 1;
defparam ram_block1a10.port_b_byte_size = 1;
defparam ram_block1a10.port_b_data_in_clock = "clock0";
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 8191;
defparam ram_block1a10.port_b_logical_ram_depth = 8192;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.port_b_write_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";
defparam ram_block1a10.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a10.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a10.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a10.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneive_ram_block ram_block1a9(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[9]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "nios_mcu_onchip_ram.hex";
defparam ram_block1a9.init_file_layout = "port_a";
defparam ram_block1a9.logical_ram_name = "nios_mcu_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_h232:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "bidir_dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 13;
defparam ram_block1a9.port_a_byte_enable_mask_width = 1;
defparam ram_block1a9.port_a_byte_size = 1;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 8191;
defparam ram_block1a9.port_a_logical_ram_depth = 8192;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 13;
defparam ram_block1a9.port_b_byte_enable_clock = "clock0";
defparam ram_block1a9.port_b_byte_enable_mask_width = 1;
defparam ram_block1a9.port_b_byte_size = 1;
defparam ram_block1a9.port_b_data_in_clock = "clock0";
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 8191;
defparam ram_block1a9.port_b_logical_ram_depth = 8192;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.port_b_write_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a9.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a9.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a9.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneive_ram_block ram_block1a8(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[8]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "nios_mcu_onchip_ram.hex";
defparam ram_block1a8.init_file_layout = "port_a";
defparam ram_block1a8.logical_ram_name = "nios_mcu_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_h232:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "bidir_dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 13;
defparam ram_block1a8.port_a_byte_enable_mask_width = 1;
defparam ram_block1a8.port_a_byte_size = 1;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 8191;
defparam ram_block1a8.port_a_logical_ram_depth = 8192;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 13;
defparam ram_block1a8.port_b_byte_enable_clock = "clock0";
defparam ram_block1a8.port_b_byte_enable_mask_width = 1;
defparam ram_block1a8.port_b_byte_size = 1;
defparam ram_block1a8.port_b_data_in_clock = "clock0";
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 8191;
defparam ram_block1a8.port_b_logical_ram_depth = 8192;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.port_b_write_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a8.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a8.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a8.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneive_ram_block ram_block1a7(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[7]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "nios_mcu_onchip_ram.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "nios_mcu_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_h232:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "bidir_dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 13;
defparam ram_block1a7.port_a_byte_enable_mask_width = 1;
defparam ram_block1a7.port_a_byte_size = 1;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 8191;
defparam ram_block1a7.port_a_logical_ram_depth = 8192;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 13;
defparam ram_block1a7.port_b_byte_enable_clock = "clock0";
defparam ram_block1a7.port_b_byte_enable_mask_width = 1;
defparam ram_block1a7.port_b_byte_size = 1;
defparam ram_block1a7.port_b_data_in_clock = "clock0";
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 8191;
defparam ram_block1a7.port_b_logical_ram_depth = 8192;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.port_b_write_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a7.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a7.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a7.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneive_ram_block ram_block1a6(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[6]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "nios_mcu_onchip_ram.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "nios_mcu_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_h232:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "bidir_dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 13;
defparam ram_block1a6.port_a_byte_enable_mask_width = 1;
defparam ram_block1a6.port_a_byte_size = 1;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 8191;
defparam ram_block1a6.port_a_logical_ram_depth = 8192;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 13;
defparam ram_block1a6.port_b_byte_enable_clock = "clock0";
defparam ram_block1a6.port_b_byte_enable_mask_width = 1;
defparam ram_block1a6.port_b_byte_size = 1;
defparam ram_block1a6.port_b_data_in_clock = "clock0";
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 8191;
defparam ram_block1a6.port_b_logical_ram_depth = 8192;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.port_b_write_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a6.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a6.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a6.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneive_ram_block ram_block1a21(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[21]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a21_PORTADATAOUT_bus),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus));
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk0_input_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.init_file = "nios_mcu_onchip_ram.hex";
defparam ram_block1a21.init_file_layout = "port_a";
defparam ram_block1a21.logical_ram_name = "nios_mcu_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_h232:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "bidir_dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 13;
defparam ram_block1a21.port_a_byte_enable_mask_width = 1;
defparam ram_block1a21.port_a_byte_size = 1;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 8191;
defparam ram_block1a21.port_a_logical_ram_depth = 8192;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock0";
defparam ram_block1a21.port_b_address_width = 13;
defparam ram_block1a21.port_b_byte_enable_clock = "clock0";
defparam ram_block1a21.port_b_byte_enable_mask_width = 1;
defparam ram_block1a21.port_b_byte_size = 1;
defparam ram_block1a21.port_b_data_in_clock = "clock0";
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 8191;
defparam ram_block1a21.port_b_logical_ram_depth = 8192;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock0";
defparam ram_block1a21.port_b_write_enable_clock = "clock0";
defparam ram_block1a21.ram_block_type = "auto";
defparam ram_block1a21.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a21.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a21.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a21.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneive_ram_block ram_block1a19(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[19]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a19_PORTADATAOUT_bus),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.init_file = "nios_mcu_onchip_ram.hex";
defparam ram_block1a19.init_file_layout = "port_a";
defparam ram_block1a19.logical_ram_name = "nios_mcu_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_h232:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "bidir_dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 13;
defparam ram_block1a19.port_a_byte_enable_mask_width = 1;
defparam ram_block1a19.port_a_byte_size = 1;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 8191;
defparam ram_block1a19.port_a_logical_ram_depth = 8192;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock0";
defparam ram_block1a19.port_b_address_width = 13;
defparam ram_block1a19.port_b_byte_enable_clock = "clock0";
defparam ram_block1a19.port_b_byte_enable_mask_width = 1;
defparam ram_block1a19.port_b_byte_size = 1;
defparam ram_block1a19.port_b_data_in_clock = "clock0";
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 8191;
defparam ram_block1a19.port_b_logical_ram_depth = 8192;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock0";
defparam ram_block1a19.port_b_write_enable_clock = "clock0";
defparam ram_block1a19.ram_block_type = "auto";
defparam ram_block1a19.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a19.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a19.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a19.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneive_ram_block ram_block1a20(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[20]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a20_PORTADATAOUT_bus),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus));
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk0_input_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.init_file = "nios_mcu_onchip_ram.hex";
defparam ram_block1a20.init_file_layout = "port_a";
defparam ram_block1a20.logical_ram_name = "nios_mcu_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_h232:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "bidir_dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 13;
defparam ram_block1a20.port_a_byte_enable_mask_width = 1;
defparam ram_block1a20.port_a_byte_size = 1;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 8191;
defparam ram_block1a20.port_a_logical_ram_depth = 8192;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock0";
defparam ram_block1a20.port_b_address_width = 13;
defparam ram_block1a20.port_b_byte_enable_clock = "clock0";
defparam ram_block1a20.port_b_byte_enable_mask_width = 1;
defparam ram_block1a20.port_b_byte_size = 1;
defparam ram_block1a20.port_b_data_in_clock = "clock0";
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 8191;
defparam ram_block1a20.port_b_logical_ram_depth = 8192;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock0";
defparam ram_block1a20.port_b_write_enable_clock = "clock0";
defparam ram_block1a20.ram_block_type = "auto";
defparam ram_block1a20.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a20.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a20.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a20.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneive_ram_block ram_block1a27(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[27]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a27_PORTADATAOUT_bus),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus));
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk0_input_clock_enable = "ena0";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.init_file = "nios_mcu_onchip_ram.hex";
defparam ram_block1a27.init_file_layout = "port_a";
defparam ram_block1a27.logical_ram_name = "nios_mcu_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_h232:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "bidir_dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 13;
defparam ram_block1a27.port_a_byte_enable_mask_width = 1;
defparam ram_block1a27.port_a_byte_size = 1;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 8191;
defparam ram_block1a27.port_a_logical_ram_depth = 8192;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock0";
defparam ram_block1a27.port_b_address_width = 13;
defparam ram_block1a27.port_b_byte_enable_clock = "clock0";
defparam ram_block1a27.port_b_byte_enable_mask_width = 1;
defparam ram_block1a27.port_b_byte_size = 1;
defparam ram_block1a27.port_b_data_in_clock = "clock0";
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 8191;
defparam ram_block1a27.port_b_logical_ram_depth = 8192;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock0";
defparam ram_block1a27.port_b_write_enable_clock = "clock0";
defparam ram_block1a27.ram_block_type = "auto";
defparam ram_block1a27.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a27.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a27.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a27.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneive_ram_block ram_block1a28(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[28]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a28_PORTADATAOUT_bus),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus));
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.clk0_input_clock_enable = "ena0";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.init_file = "nios_mcu_onchip_ram.hex";
defparam ram_block1a28.init_file_layout = "port_a";
defparam ram_block1a28.logical_ram_name = "nios_mcu_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_h232:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "bidir_dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 13;
defparam ram_block1a28.port_a_byte_enable_mask_width = 1;
defparam ram_block1a28.port_a_byte_size = 1;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 8191;
defparam ram_block1a28.port_a_logical_ram_depth = 8192;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock0";
defparam ram_block1a28.port_b_address_width = 13;
defparam ram_block1a28.port_b_byte_enable_clock = "clock0";
defparam ram_block1a28.port_b_byte_enable_mask_width = 1;
defparam ram_block1a28.port_b_byte_size = 1;
defparam ram_block1a28.port_b_data_in_clock = "clock0";
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 8191;
defparam ram_block1a28.port_b_logical_ram_depth = 8192;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock0";
defparam ram_block1a28.port_b_write_enable_clock = "clock0";
defparam ram_block1a28.ram_block_type = "auto";
defparam ram_block1a28.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a28.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a28.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a28.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneive_ram_block ram_block1a29(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[29]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a29_PORTADATAOUT_bus),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus));
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.clk0_input_clock_enable = "ena0";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.init_file = "nios_mcu_onchip_ram.hex";
defparam ram_block1a29.init_file_layout = "port_a";
defparam ram_block1a29.logical_ram_name = "nios_mcu_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_h232:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "bidir_dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 13;
defparam ram_block1a29.port_a_byte_enable_mask_width = 1;
defparam ram_block1a29.port_a_byte_size = 1;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 8191;
defparam ram_block1a29.port_a_logical_ram_depth = 8192;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock0";
defparam ram_block1a29.port_b_address_width = 13;
defparam ram_block1a29.port_b_byte_enable_clock = "clock0";
defparam ram_block1a29.port_b_byte_enable_mask_width = 1;
defparam ram_block1a29.port_b_byte_size = 1;
defparam ram_block1a29.port_b_data_in_clock = "clock0";
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 8191;
defparam ram_block1a29.port_b_logical_ram_depth = 8192;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock0";
defparam ram_block1a29.port_b_write_enable_clock = "clock0";
defparam ram_block1a29.ram_block_type = "auto";
defparam ram_block1a29.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a29.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a29.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a29.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneive_ram_block ram_block1a30(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[30]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a30_PORTADATAOUT_bus),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus));
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.clk0_input_clock_enable = "ena0";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.init_file = "nios_mcu_onchip_ram.hex";
defparam ram_block1a30.init_file_layout = "port_a";
defparam ram_block1a30.logical_ram_name = "nios_mcu_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_h232:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "bidir_dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 13;
defparam ram_block1a30.port_a_byte_enable_mask_width = 1;
defparam ram_block1a30.port_a_byte_size = 1;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 8191;
defparam ram_block1a30.port_a_logical_ram_depth = 8192;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock0";
defparam ram_block1a30.port_b_address_width = 13;
defparam ram_block1a30.port_b_byte_enable_clock = "clock0";
defparam ram_block1a30.port_b_byte_enable_mask_width = 1;
defparam ram_block1a30.port_b_byte_size = 1;
defparam ram_block1a30.port_b_data_in_clock = "clock0";
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 8191;
defparam ram_block1a30.port_b_logical_ram_depth = 8192;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock0";
defparam ram_block1a30.port_b_write_enable_clock = "clock0";
defparam ram_block1a30.ram_block_type = "auto";
defparam ram_block1a30.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a30.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a30.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a30.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneive_ram_block ram_block1a31(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(wren_b),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[31]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a31_PORTADATAOUT_bus),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus));
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.clk0_input_clock_enable = "ena0";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.init_file = "nios_mcu_onchip_ram.hex";
defparam ram_block1a31.init_file_layout = "port_a";
defparam ram_block1a31.logical_ram_name = "nios_mcu_onchip_ram:onchip_ram|altsyncram:the_altsyncram|altsyncram_h232:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "bidir_dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 13;
defparam ram_block1a31.port_a_byte_enable_mask_width = 1;
defparam ram_block1a31.port_a_byte_size = 1;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 8191;
defparam ram_block1a31.port_a_logical_ram_depth = 8192;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock0";
defparam ram_block1a31.port_b_address_width = 13;
defparam ram_block1a31.port_b_byte_enable_clock = "clock0";
defparam ram_block1a31.port_b_byte_enable_mask_width = 1;
defparam ram_block1a31.port_b_byte_size = 1;
defparam ram_block1a31.port_b_data_in_clock = "clock0";
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 8191;
defparam ram_block1a31.port_b_logical_ram_depth = 8192;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock0";
defparam ram_block1a31.port_b_write_enable_clock = "clock0";
defparam ram_block1a31.ram_block_type = "auto";
defparam ram_block1a31.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a31.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a31.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a31.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

endmodule

module nios_mcu_nios_mcu_pio_0 (
	W_alu_result_4,
	W_alu_result_3,
	W_alu_result_2,
	data_out_0,
	data_out_1,
	data_out_2,
	data_out_3,
	data_out_4,
	data_out_5,
	data_out_6,
	data_out_7,
	writedata,
	reset_n,
	Equal1,
	rst1,
	mem_used_1,
	always0,
	d_write,
	write_accepted,
	wait_latency_counter_1,
	wait_latency_counter_0,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	readdata_6,
	readdata_7,
	clk)/* synthesis synthesis_greybox=1 */;
input 	W_alu_result_4;
input 	W_alu_result_3;
input 	W_alu_result_2;
output 	data_out_0;
output 	data_out_1;
output 	data_out_2;
output 	data_out_3;
output 	data_out_4;
output 	data_out_5;
output 	data_out_6;
output 	data_out_7;
input 	[31:0] writedata;
input 	reset_n;
input 	Equal1;
input 	rst1;
input 	mem_used_1;
output 	always0;
input 	d_write;
input 	write_accepted;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_5;
output 	readdata_6;
output 	readdata_7;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~1_combout ;
wire \always0~2_combout ;


dffeas \data_out[0] (
	.clk(clk),
	.d(writedata[0]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_0),
	.prn(vcc));
defparam \data_out[0] .is_wysiwyg = "true";
defparam \data_out[0] .power_up = "low";

dffeas \data_out[1] (
	.clk(clk),
	.d(writedata[1]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_1),
	.prn(vcc));
defparam \data_out[1] .is_wysiwyg = "true";
defparam \data_out[1] .power_up = "low";

dffeas \data_out[2] (
	.clk(clk),
	.d(writedata[2]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_2),
	.prn(vcc));
defparam \data_out[2] .is_wysiwyg = "true";
defparam \data_out[2] .power_up = "low";

dffeas \data_out[3] (
	.clk(clk),
	.d(writedata[3]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_3),
	.prn(vcc));
defparam \data_out[3] .is_wysiwyg = "true";
defparam \data_out[3] .power_up = "low";

dffeas \data_out[4] (
	.clk(clk),
	.d(writedata[4]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_4),
	.prn(vcc));
defparam \data_out[4] .is_wysiwyg = "true";
defparam \data_out[4] .power_up = "low";

dffeas \data_out[5] (
	.clk(clk),
	.d(writedata[5]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_5),
	.prn(vcc));
defparam \data_out[5] .is_wysiwyg = "true";
defparam \data_out[5] .power_up = "low";

dffeas \data_out[6] (
	.clk(clk),
	.d(writedata[6]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_6),
	.prn(vcc));
defparam \data_out[6] .is_wysiwyg = "true";
defparam \data_out[6] .power_up = "low";

dffeas \data_out[7] (
	.clk(clk),
	.d(writedata[7]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~2_combout ),
	.q(data_out_7),
	.prn(vcc));
defparam \data_out[7] .is_wysiwyg = "true";
defparam \data_out[7] .power_up = "low";

cycloneive_lcell_comb \always0~0 (
	.dataa(Equal1),
	.datab(rst1),
	.datac(W_alu_result_4),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(always0),
	.cout());
defparam \always0~0 .lut_mask = 16'hEFFF;
defparam \always0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[0] (
	.dataa(data_out_0),
	.datab(gnd),
	.datac(W_alu_result_3),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(readdata_0),
	.cout());
defparam \readdata[0] .lut_mask = 16'hAFFF;
defparam \readdata[0] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[1] (
	.dataa(data_out_1),
	.datab(gnd),
	.datac(W_alu_result_3),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(readdata_1),
	.cout());
defparam \readdata[1] .lut_mask = 16'hAFFF;
defparam \readdata[1] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[2] (
	.dataa(data_out_2),
	.datab(gnd),
	.datac(W_alu_result_3),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(readdata_2),
	.cout());
defparam \readdata[2] .lut_mask = 16'hAFFF;
defparam \readdata[2] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[3] (
	.dataa(data_out_3),
	.datab(gnd),
	.datac(W_alu_result_3),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(readdata_3),
	.cout());
defparam \readdata[3] .lut_mask = 16'hAFFF;
defparam \readdata[3] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[4] (
	.dataa(data_out_4),
	.datab(gnd),
	.datac(W_alu_result_3),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(readdata_4),
	.cout());
defparam \readdata[4] .lut_mask = 16'hAFFF;
defparam \readdata[4] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[5] (
	.dataa(data_out_5),
	.datab(gnd),
	.datac(W_alu_result_3),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(readdata_5),
	.cout());
defparam \readdata[5] .lut_mask = 16'hAFFF;
defparam \readdata[5] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[6] (
	.dataa(data_out_6),
	.datab(gnd),
	.datac(W_alu_result_3),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(readdata_6),
	.cout());
defparam \readdata[6] .lut_mask = 16'hAFFF;
defparam \readdata[6] .sum_lutc_input = "datac";

cycloneive_lcell_comb \readdata[7] (
	.dataa(data_out_7),
	.datab(gnd),
	.datac(W_alu_result_3),
	.datad(W_alu_result_2),
	.cin(gnd),
	.combout(readdata_7),
	.cout());
defparam \readdata[7] .lut_mask = 16'hAFFF;
defparam \readdata[7] .sum_lutc_input = "datac";

cycloneive_lcell_comb \always0~1 (
	.dataa(d_write),
	.datab(W_alu_result_3),
	.datac(W_alu_result_2),
	.datad(write_accepted),
	.cin(gnd),
	.combout(\always0~1_combout ),
	.cout());
defparam \always0~1 .lut_mask = 16'hBFFF;
defparam \always0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always0~2 (
	.dataa(always0),
	.datab(\always0~1_combout ),
	.datac(wait_latency_counter_1),
	.datad(wait_latency_counter_0),
	.cin(gnd),
	.combout(\always0~2_combout ),
	.cout());
defparam \always0~2 .lut_mask = 16'hEFFF;
defparam \always0~2 .sum_lutc_input = "datac";

endmodule
